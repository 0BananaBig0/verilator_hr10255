module typical_example();
endmodule

