module top(A,B,ci,cco,co,SUM);
   input [23:0]A;
   input [23:0]B;
   input ci;
   inout cco;
   output co;
   output [29:0]SUM;
   wire [9:0]C;
   wire [12:0]con;
   wire [3:0]con0;
   wire [3:0]con1;
   wire [3:0]con2;
   wire [3:0]con3;
   wire cci;
   wire ccco;
   wire cc;
   wire [63:0]slongv;
   wire [127:0]longv;
   wire [255:0]llongv;
   wire zn;
   wire xn;
   wire [2:0]U1_C;
   wire U1_c_no_defined;
   wire [4:0]U1_U0_C;
   wire U1_U0_d;
   wire U1_U0_U0_d;
   wire \U1_U0_U0_U1_n_0[0] ;
   wire \U1_U0_U0_U1_n_0[1] ;
   wire \U1_U0_U0_U1_n_0[2] ;
   wire U1_U0_U0_U1_d;
   wire [15:0]\U1_U0_U0_U0_DC_output[2] ;
   wire [15:0]\U1_U0_U0_U0_DC_output[1] ;
   wire U1_U0_U1_d;
   wire \U1_U0_U1_U1_n_0[0] ;
   wire \U1_U0_U1_U1_n_0[1] ;
   wire \U1_U0_U1_U1_n_0[2] ;
   wire U1_U0_U1_U1_d;
   wire [15:0]\U1_U0_U1_U0_DC_output[2] ;
   wire [15:0]\U1_U0_U1_U0_DC_output[1] ;
   wire U1_U0_U2_d;
   wire \U1_U0_U2_U1_n_0[0] ;
   wire \U1_U0_U2_U1_n_0[1] ;
   wire \U1_U0_U2_U1_n_0[2] ;
   wire U1_U0_U2_U1_d;
   wire [15:0]\U1_U0_U2_U0_DC_output[2] ;
   wire [15:0]\U1_U0_U2_U0_DC_output[1] ;
   wire U1_U0_U3_d;
   wire \U1_U0_U3_U1_n_0[0] ;
   wire \U1_U0_U3_U1_n_0[1] ;
   wire \U1_U0_U3_U1_n_0[2] ;
   wire U1_U0_U3_U1_d;
   wire [15:0]\U1_U0_U3_U0_DC_output[2] ;
   wire [15:0]\U1_U0_U3_U0_DC_output[1] ;
   wire [4:0]U1_U1_C;
   wire U1_U1_d;
   wire U1_U1_U0_d;
   wire \U1_U1_U0_U1_n_0[0] ;
   wire \U1_U1_U0_U1_n_0[1] ;
   wire \U1_U1_U0_U1_n_0[2] ;
   wire U1_U1_U0_U1_d;
   wire [15:0]\U1_U1_U0_U0_DC_output[2] ;
   wire [15:0]\U1_U1_U0_U0_DC_output[1] ;
   wire U1_U1_U1_d;
   wire \U1_U1_U1_U1_n_0[0] ;
   wire \U1_U1_U1_U1_n_0[1] ;
   wire \U1_U1_U1_U1_n_0[2] ;
   wire U1_U1_U1_U1_d;
   wire [15:0]\U1_U1_U1_U0_DC_output[2] ;
   wire [15:0]\U1_U1_U1_U0_DC_output[1] ;
   wire U1_U1_U2_d;
   wire \U1_U1_U2_U1_n_0[0] ;
   wire \U1_U1_U2_U1_n_0[1] ;
   wire \U1_U1_U2_U1_n_0[2] ;
   wire U1_U1_U2_U1_d;
   wire [15:0]\U1_U1_U2_U0_DC_output[2] ;
   wire [15:0]\U1_U1_U2_U0_DC_output[1] ;
   wire U1_U1_U3_d;
   wire \U1_U1_U3_U1_n_0[0] ;
   wire \U1_U1_U3_U1_n_0[1] ;
   wire \U1_U1_U3_U1_n_0[2] ;
   wire U1_U1_U3_U1_d;
   wire [15:0]\U1_U1_U3_U0_DC_output[2] ;
   wire [15:0]\U1_U1_U3_U0_DC_output[1] ;
   wire [4:0]U1_U2_C;
   wire U1_U2_d;
   wire U1_U2_U0_d;
   wire \U1_U2_U0_U1_n_0[0] ;
   wire \U1_U2_U0_U1_n_0[1] ;
   wire \U1_U2_U0_U1_n_0[2] ;
   wire U1_U2_U0_U1_d;
   wire [15:0]\U1_U2_U0_U0_DC_output[2] ;
   wire [15:0]\U1_U2_U0_U0_DC_output[1] ;
   wire U1_U2_U1_d;
   wire \U1_U2_U1_U1_n_0[0] ;
   wire \U1_U2_U1_U1_n_0[1] ;
   wire \U1_U2_U1_U1_n_0[2] ;
   wire U1_U2_U1_U1_d;
   wire [15:0]\U1_U2_U1_U0_DC_output[2] ;
   wire [15:0]\U1_U2_U1_U0_DC_output[1] ;
   wire U1_U2_U2_d;
   wire \U1_U2_U2_U1_n_0[0] ;
   wire \U1_U2_U2_U1_n_0[1] ;
   wire \U1_U2_U2_U1_n_0[2] ;
   wire U1_U2_U2_U1_d;
   wire [15:0]\U1_U2_U2_U0_DC_output[2] ;
   wire [15:0]\U1_U2_U2_U0_DC_output[1] ;
   wire U1_U2_U3_d;
   wire \U1_U2_U3_U1_n_0[0] ;
   wire \U1_U2_U3_U1_n_0[1] ;
   wire \U1_U2_U3_U1_n_0[2] ;
   wire U1_U2_U3_U1_d;
   wire [15:0]\U1_U2_U3_U0_DC_output[2] ;
   wire [15:0]\U1_U2_U3_U0_DC_output[1] ;
   wire [2:0]U2_C;
   wire U2_c_no_defined;
   wire [4:0]U2_U0_C;
   wire U2_U0_d;
   wire U2_U0_U0_d;
   wire \U2_U0_U0_U1_n_0[0] ;
   wire \U2_U0_U0_U1_n_0[1] ;
   wire \U2_U0_U0_U1_n_0[2] ;
   wire U2_U0_U0_U1_d;
   wire [15:0]\U2_U0_U0_U0_DC_output[2] ;
   wire [15:0]\U2_U0_U0_U0_DC_output[1] ;
   wire U2_U0_U1_d;
   wire \U2_U0_U1_U1_n_0[0] ;
   wire \U2_U0_U1_U1_n_0[1] ;
   wire \U2_U0_U1_U1_n_0[2] ;
   wire U2_U0_U1_U1_d;
   wire [15:0]\U2_U0_U1_U0_DC_output[2] ;
   wire [15:0]\U2_U0_U1_U0_DC_output[1] ;
   wire U2_U0_U2_d;
   wire \U2_U0_U2_U1_n_0[0] ;
   wire \U2_U0_U2_U1_n_0[1] ;
   wire \U2_U0_U2_U1_n_0[2] ;
   wire U2_U0_U2_U1_d;
   wire [15:0]\U2_U0_U2_U0_DC_output[2] ;
   wire [15:0]\U2_U0_U2_U0_DC_output[1] ;
   wire U2_U0_U3_d;
   wire \U2_U0_U3_U1_n_0[0] ;
   wire \U2_U0_U3_U1_n_0[1] ;
   wire \U2_U0_U3_U1_n_0[2] ;
   wire U2_U0_U3_U1_d;
   wire [15:0]\U2_U0_U3_U0_DC_output[2] ;
   wire [15:0]\U2_U0_U3_U0_DC_output[1] ;
   wire [4:0]U2_U1_C;
   wire U2_U1_d;
   wire U2_U1_U0_d;
   wire \U2_U1_U0_U1_n_0[0] ;
   wire \U2_U1_U0_U1_n_0[1] ;
   wire \U2_U1_U0_U1_n_0[2] ;
   wire U2_U1_U0_U1_d;
   wire [15:0]\U2_U1_U0_U0_DC_output[2] ;
   wire [15:0]\U2_U1_U0_U0_DC_output[1] ;
   wire U2_U1_U1_d;
   wire \U2_U1_U1_U1_n_0[0] ;
   wire \U2_U1_U1_U1_n_0[1] ;
   wire \U2_U1_U1_U1_n_0[2] ;
   wire U2_U1_U1_U1_d;
   wire [15:0]\U2_U1_U1_U0_DC_output[2] ;
   wire [15:0]\U2_U1_U1_U0_DC_output[1] ;
   wire U2_U1_U2_d;
   wire \U2_U1_U2_U1_n_0[0] ;
   wire \U2_U1_U2_U1_n_0[1] ;
   wire \U2_U1_U2_U1_n_0[2] ;
   wire U2_U1_U2_U1_d;
   wire [15:0]\U2_U1_U2_U0_DC_output[2] ;
   wire [15:0]\U2_U1_U2_U0_DC_output[1] ;
   wire U2_U1_U3_d;
   wire \U2_U1_U3_U1_n_0[0] ;
   wire \U2_U1_U3_U1_n_0[1] ;
   wire \U2_U1_U3_U1_n_0[2] ;
   wire U2_U1_U3_U1_d;
   wire [15:0]\U2_U1_U3_U0_DC_output[2] ;
   wire [15:0]\U2_U1_U3_U0_DC_output[1] ;
   wire [4:0]U2_U2_C;
   wire U2_U2_d;
   wire U2_U2_U0_d;
   wire \U2_U2_U0_U1_n_0[0] ;
   wire \U2_U2_U0_U1_n_0[1] ;
   wire \U2_U2_U0_U1_n_0[2] ;
   wire U2_U2_U0_U1_d;
   wire [15:0]\U2_U2_U0_U0_DC_output[2] ;
   wire [15:0]\U2_U2_U0_U0_DC_output[1] ;
   wire U2_U2_U1_d;
   wire \U2_U2_U1_U1_n_0[0] ;
   wire \U2_U2_U1_U1_n_0[1] ;
   wire \U2_U2_U1_U1_n_0[2] ;
   wire U2_U2_U1_U1_d;
   wire [15:0]\U2_U2_U1_U0_DC_output[2] ;
   wire [15:0]\U2_U2_U1_U0_DC_output[1] ;
   wire U2_U2_U2_d;
   wire \U2_U2_U2_U1_n_0[0] ;
   wire \U2_U2_U2_U1_n_0[1] ;
   wire \U2_U2_U2_U1_n_0[2] ;
   wire U2_U2_U2_U1_d;
   wire [15:0]\U2_U2_U2_U0_DC_output[2] ;
   wire [15:0]\U2_U2_U2_U0_DC_output[1] ;
   wire U2_U2_U3_d;
   wire \U2_U2_U3_U1_n_0[0] ;
   wire \U2_U2_U3_U1_n_0[1] ;
   wire \U2_U2_U3_U1_n_0[2] ;
   wire U2_U2_U3_U1_d;
   wire [15:0]\U2_U2_U3_U0_DC_output[2] ;
   wire [15:0]\U2_U2_U3_U0_DC_output[1] ;
   wire U3_d;
   wire \U3_U1_n_0[0] ;
   wire \U3_U1_n_0[1] ;
   wire \U3_U1_n_0[2] ;
   wire U3_U1_d;
   wire [15:0]\U3_U0_DC_output[2] ;
   wire [15:0]\U3_U0_DC_output[1] ;
   wire U4_d;
   wire \U4_U1_n_0[0] ;
   wire \U4_U1_n_0[1] ;
   wire \U4_U1_n_0[2] ;
   wire U4_U1_d;
   wire [15:0]\U4_U0_DC_output[2] ;
   wire [15:0]\U4_U0_DC_output[1] ;
   wire \U5_n_0[0] ;
   wire \U5_n_0[1] ;
   wire \U5_n_0[2] ;
   wire U5_d;
   wire [4:0]U6_C;
   wire U6_d;
   wire U6_U0_d;
   wire \U6_U0_U1_n_0[0] ;
   wire \U6_U0_U1_n_0[1] ;
   wire \U6_U0_U1_n_0[2] ;
   wire U6_U0_U1_d;
   wire [15:0]\U6_U0_U0_DC_output[2] ;
   wire [15:0]\U6_U0_U0_DC_output[1] ;
   wire U6_U1_d;
   wire \U6_U1_U1_n_0[0] ;
   wire \U6_U1_U1_n_0[1] ;
   wire \U6_U1_U1_n_0[2] ;
   wire U6_U1_U1_d;
   wire [15:0]\U6_U1_U0_DC_output[2] ;
   wire [15:0]\U6_U1_U0_DC_output[1] ;
   wire U6_U2_d;
   wire \U6_U2_U1_n_0[0] ;
   wire \U6_U2_U1_n_0[1] ;
   wire \U6_U2_U1_n_0[2] ;
   wire U6_U2_U1_d;
   wire [15:0]\U6_U2_U0_DC_output[2] ;
   wire [15:0]\U6_U2_U0_DC_output[1] ;
   wire U6_U3_d;
   wire \U6_U3_U1_n_0[0] ;
   wire \U6_U3_U1_n_0[1] ;
   wire \U6_U3_U1_n_0[2] ;
   wire U6_U3_U1_d;
   wire [15:0]\U6_U3_U0_DC_output[2] ;
   wire [15:0]\U6_U3_U0_DC_output[1] ;
   wire [4:0]U8_C;
   wire U8_d;
   wire U8_U0_d;
   wire \U8_U0_U1_n_0[0] ;
   wire \U8_U0_U1_n_0[1] ;
   wire \U8_U0_U1_n_0[2] ;
   wire U8_U0_U1_d;
   wire [15:0]\U8_U0_U0_DC_output[2] ;
   wire [15:0]\U8_U0_U0_DC_output[1] ;
   wire U8_U1_d;
   wire \U8_U1_U1_n_0[0] ;
   wire \U8_U1_U1_n_0[1] ;
   wire \U8_U1_U1_n_0[2] ;
   wire U8_U1_U1_d;
   wire [15:0]\U8_U1_U0_DC_output[2] ;
   wire [15:0]\U8_U1_U0_DC_output[1] ;
   wire U8_U2_d;
   wire \U8_U2_U1_n_0[0] ;
   wire \U8_U2_U1_n_0[1] ;
   wire \U8_U2_U1_n_0[2] ;
   wire U8_U2_U1_d;
   wire [15:0]\U8_U2_U0_DC_output[2] ;
   wire [15:0]\U8_U2_U0_DC_output[1] ;
   wire U8_U3_d;
   wire \U8_U3_U1_n_0[0] ;
   wire \U8_U3_U1_n_0[1] ;
   wire \U8_U3_U1_n_0[2] ;
   wire U8_U3_U1_d;
   wire [15:0]\U8_U3_U0_DC_output[2] ;
   wire [15:0]\U8_U3_U0_DC_output[1] ;
   wire [2:0]U9_C;
   wire U9_c_no_defined;
   wire [4:0]U9_U0_C;
   wire U9_U0_d;
   wire U9_U0_U0_d;
   wire \U9_U0_U0_U1_n_0[0] ;
   wire \U9_U0_U0_U1_n_0[1] ;
   wire \U9_U0_U0_U1_n_0[2] ;
   wire U9_U0_U0_U1_d;
   wire [15:0]\U9_U0_U0_U0_DC_output[2] ;
   wire [15:0]\U9_U0_U0_U0_DC_output[1] ;
   wire U9_U0_U1_d;
   wire \U9_U0_U1_U1_n_0[0] ;
   wire \U9_U0_U1_U1_n_0[1] ;
   wire \U9_U0_U1_U1_n_0[2] ;
   wire U9_U0_U1_U1_d;
   wire [15:0]\U9_U0_U1_U0_DC_output[2] ;
   wire [15:0]\U9_U0_U1_U0_DC_output[1] ;
   wire U9_U0_U2_d;
   wire \U9_U0_U2_U1_n_0[0] ;
   wire \U9_U0_U2_U1_n_0[1] ;
   wire \U9_U0_U2_U1_n_0[2] ;
   wire U9_U0_U2_U1_d;
   wire [15:0]\U9_U0_U2_U0_DC_output[2] ;
   wire [15:0]\U9_U0_U2_U0_DC_output[1] ;
   wire U9_U0_U3_d;
   wire \U9_U0_U3_U1_n_0[0] ;
   wire \U9_U0_U3_U1_n_0[1] ;
   wire \U9_U0_U3_U1_n_0[2] ;
   wire U9_U0_U3_U1_d;
   wire [15:0]\U9_U0_U3_U0_DC_output[2] ;
   wire [15:0]\U9_U0_U3_U0_DC_output[1] ;
   wire [4:0]U9_U1_C;
   wire U9_U1_d;
   wire U9_U1_U0_d;
   wire \U9_U1_U0_U1_n_0[0] ;
   wire \U9_U1_U0_U1_n_0[1] ;
   wire \U9_U1_U0_U1_n_0[2] ;
   wire U9_U1_U0_U1_d;
   wire [15:0]\U9_U1_U0_U0_DC_output[2] ;
   wire [15:0]\U9_U1_U0_U0_DC_output[1] ;
   wire U9_U1_U1_d;
   wire \U9_U1_U1_U1_n_0[0] ;
   wire \U9_U1_U1_U1_n_0[1] ;
   wire \U9_U1_U1_U1_n_0[2] ;
   wire U9_U1_U1_U1_d;
   wire [15:0]\U9_U1_U1_U0_DC_output[2] ;
   wire [15:0]\U9_U1_U1_U0_DC_output[1] ;
   wire U9_U1_U2_d;
   wire \U9_U1_U2_U1_n_0[0] ;
   wire \U9_U1_U2_U1_n_0[1] ;
   wire \U9_U1_U2_U1_n_0[2] ;
   wire U9_U1_U2_U1_d;
   wire [15:0]\U9_U1_U2_U0_DC_output[2] ;
   wire [15:0]\U9_U1_U2_U0_DC_output[1] ;
   wire U9_U1_U3_d;
   wire \U9_U1_U3_U1_n_0[0] ;
   wire \U9_U1_U3_U1_n_0[1] ;
   wire \U9_U1_U3_U1_n_0[2] ;
   wire U9_U1_U3_U1_d;
   wire [15:0]\U9_U1_U3_U0_DC_output[2] ;
   wire [15:0]\U9_U1_U3_U0_DC_output[1] ;
   wire [4:0]U9_U2_C;
   wire U9_U2_d;
   wire U9_U2_U0_d;
   wire \U9_U2_U0_U1_n_0[0] ;
   wire \U9_U2_U0_U1_n_0[1] ;
   wire \U9_U2_U0_U1_n_0[2] ;
   wire U9_U2_U0_U1_d;
   wire [15:0]\U9_U2_U0_U0_DC_output[2] ;
   wire [15:0]\U9_U2_U0_U0_DC_output[1] ;
   wire U9_U2_U1_d;
   wire \U9_U2_U1_U1_n_0[0] ;
   wire \U9_U2_U1_U1_n_0[1] ;
   wire \U9_U2_U1_U1_n_0[2] ;
   wire U9_U2_U1_U1_d;
   wire [15:0]\U9_U2_U1_U0_DC_output[2] ;
   wire [15:0]\U9_U2_U1_U0_DC_output[1] ;
   wire U9_U2_U2_d;
   wire \U9_U2_U2_U1_n_0[0] ;
   wire \U9_U2_U2_U1_n_0[1] ;
   wire \U9_U2_U2_U1_n_0[2] ;
   wire U9_U2_U2_U1_d;
   wire [15:0]\U9_U2_U2_U0_DC_output[2] ;
   wire [15:0]\U9_U2_U2_U0_DC_output[1] ;
   wire U9_U2_U3_d;
   wire \U9_U2_U3_U1_n_0[0] ;
   wire \U9_U2_U3_U1_n_0[1] ;
   wire \U9_U2_U3_U1_n_0[2] ;
   wire U9_U2_U3_U1_d;
   wire [15:0]\U9_U2_U3_U0_DC_output[2] ;
   wire [15:0]\U9_U2_U3_U0_DC_output[1] ;
  assign C[0] = 1'b0;
  assign C[2] = 1'b1;
  assign C[3] = ci;
  assign C[4] = 1'b0;
  assign co = C[6];
  assign cci = ci;
  assign ccco = C[5];
  assign cco = ccco;
  assign con[0] = cci;
  assign con[1] = 1'b1;
  assign con[2] = 1'b1;
  assign con[3] = cco;
  assign con[4] = 1'b0;
  assign con[5] = ci;
  assign con[9] = 1'b0;
  assign con[8] = 1'b0;
  assign con[7] = 1'b1;
  assign con[6] = 1'b1;
  assign con[10] = 1'b0;
  assign con[11] = 1'b0;
  assign con[12] = 1'b1;
  assign con0[0] = 1'b0;
  assign con0[3] = 1'b1;
  assign con0[1] = 1'b1;
  assign con0[2] = cco;
  assign con1[0] = 1'b0;
  assign con1[1] = 1'b0;
  assign con1[3] = 1'b1;
  assign con1[2] = cco;
  assign con2[0] = 1'b0;
  assign con2[1] = 1'b0;
  assign con2[2] = cco;
  assign con2[3] = 1'b1;
  assign con3[3] = 1'b1;
  assign con3[2] = con[8];
  assign con3[1] = con[7];
  assign con3[0] = con[6];
  assign zn = 1'bz;
  assign xn = 1'bx;
  assign cc = 1'b1;
  assign slongv[63] = 1'b0;
  assign slongv[62] = 1'b0;
  assign slongv[61] = 1'b0;
  assign slongv[60] = 1'b0;
  assign slongv[59] = 1'b0;
  assign slongv[58] = 1'b0;
  assign slongv[57] = 1'b0;
  assign slongv[56] = 1'b0;
  assign slongv[55] = 1'b0;
  assign slongv[54] = 1'b0;
  assign slongv[53] = 1'b0;
  assign slongv[52] = 1'b0;
  assign slongv[51] = 1'b0;
  assign slongv[50] = 1'b0;
  assign slongv[49] = 1'b0;
  assign slongv[48] = 1'b0;
  assign slongv[47] = 1'b0;
  assign slongv[46] = 1'b0;
  assign slongv[45] = 1'b0;
  assign slongv[44] = 1'b0;
  assign slongv[43] = 1'b0;
  assign slongv[42] = 1'b0;
  assign slongv[41] = 1'b0;
  assign slongv[40] = 1'b0;
  assign slongv[39] = 1'b0;
  assign slongv[38] = 1'b0;
  assign slongv[37] = 1'b0;
  assign slongv[36] = 1'b0;
  assign slongv[35] = 1'b0;
  assign slongv[34] = 1'b0;
  assign slongv[33] = 1'b1;
  assign slongv[32] = 1'b0;
  assign slongv[31] = 1'b0;
  assign slongv[30] = 1'b0;
  assign slongv[29] = 1'b0;
  assign slongv[28] = 1'b0;
  assign slongv[27] = 1'b0;
  assign slongv[26] = 1'b0;
  assign slongv[25] = 1'b0;
  assign slongv[24] = 1'b0;
  assign slongv[23] = 1'b0;
  assign slongv[22] = 1'b0;
  assign slongv[21] = 1'b0;
  assign slongv[20] = 1'b0;
  assign slongv[19] = 1'b0;
  assign slongv[18] = 1'b0;
  assign slongv[17] = 1'b0;
  assign slongv[16] = 1'b0;
  assign slongv[15] = 1'b0;
  assign slongv[14] = 1'b0;
  assign slongv[13] = 1'b0;
  assign slongv[12] = 1'b0;
  assign slongv[11] = 1'b0;
  assign slongv[10] = 1'b0;
  assign slongv[9] = 1'b0;
  assign slongv[8] = 1'b0;
  assign slongv[7] = 1'b0;
  assign slongv[6] = 1'b0;
  assign slongv[5] = 1'b0;
  assign slongv[4] = 1'b0;
  assign slongv[3] = 1'b0;
  assign slongv[2] = 1'b0;
  assign slongv[1] = 1'b0;
  assign slongv[0] = 1'b1;
  assign longv[127] = 1'b0;
  assign longv[126] = 1'b0;
  assign longv[125] = 1'b0;
  assign longv[124] = 1'b0;
  assign longv[123] = 1'b0;
  assign longv[122] = 1'b0;
  assign longv[121] = 1'b0;
  assign longv[120] = 1'b0;
  assign longv[119] = 1'b0;
  assign longv[118] = 1'b0;
  assign longv[117] = 1'b0;
  assign longv[116] = 1'b0;
  assign longv[115] = 1'b0;
  assign longv[114] = 1'b0;
  assign longv[113] = 1'b0;
  assign longv[112] = 1'b0;
  assign longv[111] = 1'b0;
  assign longv[110] = 1'b0;
  assign longv[109] = 1'b0;
  assign longv[108] = 1'b0;
  assign longv[107] = 1'b0;
  assign longv[106] = 1'b0;
  assign longv[105] = 1'b0;
  assign longv[104] = 1'b0;
  assign longv[103] = 1'b0;
  assign longv[102] = 1'b0;
  assign longv[101] = 1'b0;
  assign longv[100] = 1'b0;
  assign longv[99] = 1'b0;
  assign longv[98] = 1'b0;
  assign longv[97] = 1'b1;
  assign longv[96] = 1'b0;
  assign longv[95] = 1'b0;
  assign longv[94] = 1'b0;
  assign longv[93] = 1'b0;
  assign longv[92] = 1'b0;
  assign longv[91] = 1'b0;
  assign longv[90] = 1'b0;
  assign longv[89] = 1'b0;
  assign longv[88] = 1'b0;
  assign longv[87] = 1'b0;
  assign longv[86] = 1'b0;
  assign longv[85] = 1'b0;
  assign longv[84] = 1'b0;
  assign longv[83] = 1'b0;
  assign longv[82] = 1'b0;
  assign longv[81] = 1'b0;
  assign longv[80] = 1'b0;
  assign longv[79] = 1'b0;
  assign longv[78] = 1'b0;
  assign longv[77] = 1'b0;
  assign longv[76] = 1'b0;
  assign longv[75] = 1'b0;
  assign longv[74] = 1'b0;
  assign longv[73] = 1'b0;
  assign longv[72] = 1'b0;
  assign longv[71] = 1'b0;
  assign longv[70] = 1'b0;
  assign longv[69] = 1'b0;
  assign longv[68] = 1'b0;
  assign longv[67] = 1'b0;
  assign longv[66] = 1'b0;
  assign longv[65] = 1'b1;
  assign longv[64] = 1'b0;
  assign longv[63] = 1'b0;
  assign longv[62] = 1'b0;
  assign longv[61] = 1'b0;
  assign longv[60] = 1'b0;
  assign longv[59] = 1'b0;
  assign longv[58] = 1'b0;
  assign longv[57] = 1'b0;
  assign longv[56] = 1'b0;
  assign longv[55] = 1'b0;
  assign longv[54] = 1'b0;
  assign longv[53] = 1'b0;
  assign longv[52] = 1'b0;
  assign longv[51] = 1'b0;
  assign longv[50] = 1'b0;
  assign longv[49] = 1'b0;
  assign longv[48] = 1'b0;
  assign longv[47] = 1'b0;
  assign longv[46] = 1'b0;
  assign longv[45] = 1'b0;
  assign longv[44] = 1'b0;
  assign longv[43] = 1'b0;
  assign longv[42] = 1'b0;
  assign longv[41] = 1'b0;
  assign longv[40] = 1'b0;
  assign longv[39] = 1'b0;
  assign longv[38] = 1'b0;
  assign longv[37] = 1'b0;
  assign longv[36] = 1'b0;
  assign longv[35] = 1'b0;
  assign longv[34] = 1'b0;
  assign longv[33] = 1'b1;
  assign longv[32] = 1'b0;
  assign longv[31] = 1'b0;
  assign longv[30] = 1'b0;
  assign longv[29] = 1'b0;
  assign longv[28] = 1'b0;
  assign longv[27] = 1'b0;
  assign longv[26] = 1'b0;
  assign longv[25] = 1'b0;
  assign longv[24] = 1'b0;
  assign longv[23] = 1'b0;
  assign longv[22] = 1'b0;
  assign longv[21] = 1'b0;
  assign longv[20] = 1'b0;
  assign longv[19] = 1'b0;
  assign longv[18] = 1'b0;
  assign longv[17] = 1'b0;
  assign longv[16] = 1'b0;
  assign longv[15] = 1'b0;
  assign longv[14] = 1'b0;
  assign longv[13] = 1'b0;
  assign longv[12] = 1'b0;
  assign longv[11] = 1'b0;
  assign longv[10] = 1'b0;
  assign longv[9] = 1'b0;
  assign longv[8] = 1'b0;
  assign longv[7] = 1'b0;
  assign longv[6] = 1'b0;
  assign longv[5] = 1'b0;
  assign longv[4] = 1'b0;
  assign longv[3] = 1'b0;
  assign longv[2] = 1'b0;
  assign longv[1] = 1'b0;
  assign longv[0] = 1'b1;
  assign llongv[255] = 1'b0;
  assign llongv[254] = 1'b0;
  assign llongv[253] = 1'b0;
  assign llongv[252] = 1'b0;
  assign llongv[251] = 1'b0;
  assign llongv[250] = 1'b0;
  assign llongv[249] = 1'b0;
  assign llongv[248] = 1'b0;
  assign llongv[247] = 1'b0;
  assign llongv[246] = 1'b0;
  assign llongv[245] = 1'b0;
  assign llongv[244] = 1'b0;
  assign llongv[243] = 1'b0;
  assign llongv[242] = 1'b0;
  assign llongv[241] = 1'b0;
  assign llongv[240] = 1'b0;
  assign llongv[239] = 1'b0;
  assign llongv[238] = 1'b0;
  assign llongv[237] = 1'b0;
  assign llongv[236] = 1'b0;
  assign llongv[235] = 1'b0;
  assign llongv[234] = 1'b0;
  assign llongv[233] = 1'b0;
  assign llongv[232] = 1'b0;
  assign llongv[231] = 1'b0;
  assign llongv[230] = 1'b0;
  assign llongv[229] = 1'b0;
  assign llongv[228] = 1'b0;
  assign llongv[227] = 1'b0;
  assign llongv[226] = 1'b0;
  assign llongv[225] = 1'b1;
  assign llongv[224] = 1'b0;
  assign llongv[223] = 1'b0;
  assign llongv[222] = 1'b0;
  assign llongv[221] = 1'b0;
  assign llongv[220] = 1'b0;
  assign llongv[219] = 1'b0;
  assign llongv[218] = 1'b0;
  assign llongv[217] = 1'b0;
  assign llongv[216] = 1'b0;
  assign llongv[215] = 1'b0;
  assign llongv[214] = 1'b0;
  assign llongv[213] = 1'b0;
  assign llongv[212] = 1'b0;
  assign llongv[211] = 1'b0;
  assign llongv[210] = 1'b0;
  assign llongv[209] = 1'b0;
  assign llongv[208] = 1'b0;
  assign llongv[207] = 1'b0;
  assign llongv[206] = 1'b0;
  assign llongv[205] = 1'b0;
  assign llongv[204] = 1'b0;
  assign llongv[203] = 1'b0;
  assign llongv[202] = 1'b0;
  assign llongv[201] = 1'b0;
  assign llongv[200] = 1'b0;
  assign llongv[199] = 1'b0;
  assign llongv[198] = 1'b0;
  assign llongv[197] = 1'b0;
  assign llongv[196] = 1'b0;
  assign llongv[195] = 1'b0;
  assign llongv[194] = 1'b0;
  assign llongv[193] = 1'b0;
  assign llongv[192] = 1'b1;
  assign llongv[191] = 1'b0;
  assign llongv[190] = 1'b0;
  assign llongv[189] = 1'b0;
  assign llongv[188] = 1'b0;
  assign llongv[187] = 1'b0;
  assign llongv[186] = 1'b0;
  assign llongv[185] = 1'b0;
  assign llongv[184] = 1'b0;
  assign llongv[183] = 1'b0;
  assign llongv[182] = 1'b0;
  assign llongv[181] = 1'b0;
  assign llongv[180] = 1'b0;
  assign llongv[179] = 1'b0;
  assign llongv[178] = 1'b0;
  assign llongv[177] = 1'b0;
  assign llongv[176] = 1'b0;
  assign llongv[175] = 1'b0;
  assign llongv[174] = 1'b0;
  assign llongv[173] = 1'b0;
  assign llongv[172] = 1'b0;
  assign llongv[171] = 1'b0;
  assign llongv[170] = 1'b0;
  assign llongv[169] = 1'b0;
  assign llongv[168] = 1'b0;
  assign llongv[167] = 1'b0;
  assign llongv[166] = 1'b0;
  assign llongv[165] = 1'b0;
  assign llongv[164] = 1'b0;
  assign llongv[163] = 1'b0;
  assign llongv[162] = 1'b0;
  assign llongv[161] = 1'b1;
  assign llongv[160] = 1'b0;
  assign llongv[159] = 1'b0;
  assign llongv[158] = 1'b0;
  assign llongv[157] = 1'b0;
  assign llongv[156] = 1'b0;
  assign llongv[155] = 1'b0;
  assign llongv[154] = 1'b0;
  assign llongv[153] = 1'b0;
  assign llongv[152] = 1'b0;
  assign llongv[151] = 1'b0;
  assign llongv[150] = 1'b0;
  assign llongv[149] = 1'b0;
  assign llongv[148] = 1'b0;
  assign llongv[147] = 1'b0;
  assign llongv[146] = 1'b0;
  assign llongv[145] = 1'b0;
  assign llongv[144] = 1'b0;
  assign llongv[143] = 1'b0;
  assign llongv[142] = 1'b0;
  assign llongv[141] = 1'b0;
  assign llongv[140] = 1'b0;
  assign llongv[139] = 1'b0;
  assign llongv[138] = 1'b0;
  assign llongv[137] = 1'b0;
  assign llongv[136] = 1'b0;
  assign llongv[135] = 1'b0;
  assign llongv[134] = 1'b0;
  assign llongv[133] = 1'b0;
  assign llongv[132] = 1'b0;
  assign llongv[131] = 1'b0;
  assign llongv[130] = 1'b0;
  assign llongv[129] = 1'b1;
  assign llongv[128] = 1'b0;
  assign llongv[127] = 1'b0;
  assign llongv[126] = 1'b0;
  assign llongv[125] = 1'b0;
  assign llongv[124] = 1'b0;
  assign llongv[123] = 1'b0;
  assign llongv[122] = 1'b0;
  assign llongv[121] = 1'b0;
  assign llongv[120] = 1'b0;
  assign llongv[119] = 1'b0;
  assign llongv[118] = 1'b0;
  assign llongv[117] = 1'b0;
  assign llongv[116] = 1'b0;
  assign llongv[115] = 1'b0;
  assign llongv[114] = 1'b0;
  assign llongv[113] = 1'b0;
  assign llongv[112] = 1'b0;
  assign llongv[111] = 1'b0;
  assign llongv[110] = 1'b0;
  assign llongv[109] = 1'b0;
  assign llongv[108] = 1'b0;
  assign llongv[107] = 1'b0;
  assign llongv[106] = 1'b0;
  assign llongv[105] = 1'b0;
  assign llongv[104] = 1'b0;
  assign llongv[103] = 1'b0;
  assign llongv[102] = 1'b0;
  assign llongv[101] = 1'b0;
  assign llongv[100] = 1'b0;
  assign llongv[99] = 1'b0;
  assign llongv[98] = 1'b0;
  assign llongv[97] = 1'b1;
  assign llongv[96] = 1'b0;
  assign llongv[95] = 1'b0;
  assign llongv[94] = 1'b0;
  assign llongv[93] = 1'b0;
  assign llongv[92] = 1'b0;
  assign llongv[91] = 1'b0;
  assign llongv[90] = 1'b0;
  assign llongv[89] = 1'b0;
  assign llongv[88] = 1'b0;
  assign llongv[87] = 1'b0;
  assign llongv[86] = 1'b0;
  assign llongv[85] = 1'b0;
  assign llongv[84] = 1'b0;
  assign llongv[83] = 1'b0;
  assign llongv[82] = 1'b0;
  assign llongv[81] = 1'b0;
  assign llongv[80] = 1'b0;
  assign llongv[79] = 1'b0;
  assign llongv[78] = 1'b0;
  assign llongv[77] = 1'b0;
  assign llongv[76] = 1'b0;
  assign llongv[75] = 1'b0;
  assign llongv[74] = 1'b0;
  assign llongv[73] = 1'b0;
  assign llongv[72] = 1'b0;
  assign llongv[71] = 1'b0;
  assign llongv[70] = 1'b0;
  assign llongv[69] = 1'b0;
  assign llongv[68] = 1'b0;
  assign llongv[67] = 1'b0;
  assign llongv[66] = 1'b0;
  assign llongv[65] = 1'b0;
  assign llongv[64] = 1'b1;
  assign llongv[63] = 1'b0;
  assign llongv[62] = 1'b0;
  assign llongv[61] = 1'b0;
  assign llongv[60] = 1'b0;
  assign llongv[59] = 1'b0;
  assign llongv[58] = 1'b0;
  assign llongv[57] = 1'b0;
  assign llongv[56] = 1'b0;
  assign llongv[55] = 1'b0;
  assign llongv[54] = 1'b0;
  assign llongv[53] = 1'b0;
  assign llongv[52] = 1'b0;
  assign llongv[51] = 1'b0;
  assign llongv[50] = 1'b0;
  assign llongv[49] = 1'b0;
  assign llongv[48] = 1'b0;
  assign llongv[47] = 1'b0;
  assign llongv[46] = 1'b0;
  assign llongv[45] = 1'b0;
  assign llongv[44] = 1'b0;
  assign llongv[43] = 1'b0;
  assign llongv[42] = 1'b0;
  assign llongv[41] = 1'b0;
  assign llongv[40] = 1'b0;
  assign llongv[39] = 1'b0;
  assign llongv[38] = 1'b0;
  assign llongv[37] = 1'b0;
  assign llongv[36] = 1'b0;
  assign llongv[35] = 1'b0;
  assign llongv[34] = 1'b0;
  assign llongv[33] = 1'b1;
  assign llongv[32] = 1'b0;
  assign llongv[31] = 1'b0;
  assign llongv[30] = 1'b0;
  assign llongv[29] = 1'b0;
  assign llongv[28] = 1'b0;
  assign llongv[27] = 1'b0;
  assign llongv[26] = 1'b0;
  assign llongv[25] = 1'b0;
  assign llongv[24] = 1'b0;
  assign llongv[23] = 1'b0;
  assign llongv[22] = 1'b0;
  assign llongv[21] = 1'b0;
  assign llongv[20] = 1'b0;
  assign llongv[19] = 1'b0;
  assign llongv[18] = 1'b0;
  assign llongv[17] = 1'b0;
  assign llongv[16] = 1'b0;
  assign llongv[15] = 1'b0;
  assign llongv[14] = 1'b0;
  assign llongv[13] = 1'b0;
  assign llongv[12] = 1'b0;
  assign llongv[11] = 1'b0;
  assign llongv[10] = 1'b0;
  assign llongv[9] = 1'b0;
  assign llongv[8] = 1'b0;
  assign llongv[7] = 1'b0;
  assign llongv[6] = 1'b0;
  assign llongv[5] = 1'b0;
  assign llongv[4] = 1'b0;
  assign llongv[3] = 1'b0;
  assign llongv[2] = 1'b0;
  assign llongv[1] = 1'b0;
  assign llongv[0] = 1'b1;
  assign U1_C[0] = C[9];
  assign C[5] = U1_c_no_defined;
  assign U1_U0_d = 1'b0;
  assign U1_U0_U0_d = 1'b0;
  assign U1_U0_U0_U1_d = 1'b0;
  assign \U1_U0_U0_U0_DC_output[2] [14] = 1'b0;
  assign U1_U0_U1_d = 1'b0;
  assign U1_U0_U1_U1_d = 1'b0;
  assign \U1_U0_U1_U0_DC_output[2] [14] = 1'b0;
  assign U1_U0_U2_d = 1'b0;
  assign U1_U0_U2_U1_d = 1'b0;
  assign \U1_U0_U2_U0_DC_output[2] [14] = 1'b0;
  assign U1_U0_U3_d = 1'b0;
  assign U1_U0_U3_U1_d = 1'b0;
  assign \U1_U0_U3_U0_DC_output[2] [14] = 1'b0;
  assign U1_U1_d = 1'b0;
  assign U1_U1_U0_d = 1'b0;
  assign U1_U1_U0_U1_d = 1'b0;
  assign \U1_U1_U0_U0_DC_output[2] [14] = 1'b0;
  assign U1_U1_U1_d = 1'b0;
  assign U1_U1_U1_U1_d = 1'b0;
  assign \U1_U1_U1_U0_DC_output[2] [14] = 1'b0;
  assign U1_U1_U2_d = 1'b0;
  assign U1_U1_U2_U1_d = 1'b0;
  assign \U1_U1_U2_U0_DC_output[2] [14] = 1'b0;
  assign U1_U1_U3_d = 1'b0;
  assign U1_U1_U3_U1_d = 1'b0;
  assign \U1_U1_U3_U0_DC_output[2] [14] = 1'b0;
  assign U1_U2_d = 1'b0;
  assign U1_U2_U0_d = 1'b0;
  assign U1_U2_U0_U1_d = 1'b0;
  assign \U1_U2_U0_U0_DC_output[2] [14] = 1'b0;
  assign U1_U2_U1_d = 1'b0;
  assign U1_U2_U1_U1_d = 1'b0;
  assign \U1_U2_U1_U0_DC_output[2] [14] = 1'b0;
  assign U1_U2_U2_d = 1'b0;
  assign U1_U2_U2_U1_d = 1'b0;
  assign \U1_U2_U2_U0_DC_output[2] [14] = 1'b0;
  assign U1_U2_U3_d = 1'b0;
  assign U1_U2_U3_U1_d = 1'b0;
  assign \U1_U2_U3_U0_DC_output[2] [14] = 1'b0;
  assign U2_C[0] = C[5];
  assign C[6] = U2_c_no_defined;
  assign U2_U0_d = 1'b0;
  assign U2_U0_U0_d = 1'b0;
  assign U2_U0_U0_U1_d = 1'b0;
  assign \U2_U0_U0_U0_DC_output[2] [14] = 1'b0;
  assign U2_U0_U1_d = 1'b0;
  assign U2_U0_U1_U1_d = 1'b0;
  assign \U2_U0_U1_U0_DC_output[2] [14] = 1'b0;
  assign U2_U0_U2_d = 1'b0;
  assign U2_U0_U2_U1_d = 1'b0;
  assign \U2_U0_U2_U0_DC_output[2] [14] = 1'b0;
  assign U2_U0_U3_d = 1'b0;
  assign U2_U0_U3_U1_d = 1'b0;
  assign \U2_U0_U3_U0_DC_output[2] [14] = 1'b0;
  assign U2_U1_d = 1'b0;
  assign U2_U1_U0_d = 1'b0;
  assign U2_U1_U0_U1_d = 1'b0;
  assign \U2_U1_U0_U0_DC_output[2] [14] = 1'b0;
  assign U2_U1_U1_d = 1'b0;
  assign U2_U1_U1_U1_d = 1'b0;
  assign \U2_U1_U1_U0_DC_output[2] [14] = 1'b0;
  assign U2_U1_U2_d = 1'b0;
  assign U2_U1_U2_U1_d = 1'b0;
  assign \U2_U1_U2_U0_DC_output[2] [14] = 1'b0;
  assign U2_U1_U3_d = 1'b0;
  assign U2_U1_U3_U1_d = 1'b0;
  assign \U2_U1_U3_U0_DC_output[2] [14] = 1'b0;
  assign U2_U2_d = 1'b0;
  assign U2_U2_U0_d = 1'b0;
  assign U2_U2_U0_U1_d = 1'b0;
  assign \U2_U2_U0_U0_DC_output[2] [14] = 1'b0;
  assign U2_U2_U1_d = 1'b0;
  assign U2_U2_U1_U1_d = 1'b0;
  assign \U2_U2_U1_U0_DC_output[2] [14] = 1'b0;
  assign U2_U2_U2_d = 1'b0;
  assign U2_U2_U2_U1_d = 1'b0;
  assign \U2_U2_U2_U0_DC_output[2] [14] = 1'b0;
  assign U2_U2_U3_d = 1'b0;
  assign U2_U2_U3_U1_d = 1'b0;
  assign \U2_U2_U3_U0_DC_output[2] [14] = 1'b0;
  assign U3_d = 1'b0;
  assign U3_U1_d = 1'b0;
  assign \U3_U0_DC_output[2] [14] = 1'b0;
  assign U4_d = 1'b0;
  assign U4_U1_d = 1'b0;
  assign \U4_U0_DC_output[2] [14] = 1'b0;
  assign U5_d = 1'b0;
  assign U6_d = 1'b0;
  assign U6_U0_d = 1'b0;
  assign U6_U0_U1_d = 1'b0;
  assign \U6_U0_U0_DC_output[2] [14] = 1'b0;
  assign U6_U1_d = 1'b0;
  assign U6_U1_U1_d = 1'b0;
  assign \U6_U1_U0_DC_output[2] [14] = 1'b0;
  assign U6_U2_d = 1'b0;
  assign U6_U2_U1_d = 1'b0;
  assign \U6_U2_U0_DC_output[2] [14] = 1'b0;
  assign U6_U3_d = 1'b0;
  assign U6_U3_U1_d = 1'b0;
  assign \U6_U3_U0_DC_output[2] [14] = 1'b0;
  assign U8_d = 1'b0;
  assign U8_U0_d = 1'b0;
  assign U8_U0_U1_d = 1'b0;
  assign \U8_U0_U0_DC_output[2] [14] = 1'b0;
  assign U8_U1_d = 1'b0;
  assign U8_U1_U1_d = 1'b0;
  assign \U8_U1_U0_DC_output[2] [14] = 1'b0;
  assign U8_U2_d = 1'b0;
  assign U8_U2_U1_d = 1'b0;
  assign \U8_U2_U0_DC_output[2] [14] = 1'b0;
  assign U8_U3_d = 1'b0;
  assign U8_U3_U1_d = 1'b0;
  assign \U8_U3_U0_DC_output[2] [14] = 1'b0;
  assign U9_C[0] = 1'bz;
  assign U9_U0_d = 1'b0;
  assign U9_U0_U0_d = 1'b0;
  assign U9_U0_U0_U1_d = 1'b0;
  assign \U9_U0_U0_U0_DC_output[2] [14] = 1'b0;
  assign U9_U0_U1_d = 1'b0;
  assign U9_U0_U1_U1_d = 1'b0;
  assign \U9_U0_U1_U0_DC_output[2] [14] = 1'b0;
  assign U9_U0_U2_d = 1'b0;
  assign U9_U0_U2_U1_d = 1'b0;
  assign \U9_U0_U2_U0_DC_output[2] [14] = 1'b0;
  assign U9_U0_U3_d = 1'b0;
  assign U9_U0_U3_U1_d = 1'b0;
  assign \U9_U0_U3_U0_DC_output[2] [14] = 1'b0;
  assign U9_U1_d = 1'b0;
  assign U9_U1_U0_d = 1'b0;
  assign U9_U1_U0_U1_d = 1'b0;
  assign \U9_U1_U0_U0_DC_output[2] [14] = 1'b0;
  assign U9_U1_U1_d = 1'b0;
  assign U9_U1_U1_U1_d = 1'b0;
  assign \U9_U1_U1_U0_DC_output[2] [14] = 1'b0;
  assign U9_U1_U2_d = 1'b0;
  assign U9_U1_U2_U1_d = 1'b0;
  assign \U9_U1_U2_U0_DC_output[2] [14] = 1'b0;
  assign U9_U1_U3_d = 1'b0;
  assign U9_U1_U3_U1_d = 1'b0;
  assign \U9_U1_U3_U0_DC_output[2] [14] = 1'b0;
  assign U9_U2_d = 1'b0;
  assign U9_U2_U0_d = 1'b0;
  assign U9_U2_U0_U1_d = 1'b0;
  assign \U9_U2_U0_U0_DC_output[2] [14] = 1'b0;
  assign U9_U2_U1_d = 1'b0;
  assign U9_U2_U1_U1_d = 1'b0;
  assign \U9_U2_U1_U0_DC_output[2] [14] = 1'b0;
  assign U9_U2_U2_d = 1'b0;
  assign U9_U2_U2_U1_d = 1'b0;
  assign \U9_U2_U2_U0_DC_output[2] [14] = 1'b0;
  assign U9_U2_U3_d = 1'b0;
  assign U9_U2_U3_U1_d = 1'b0;
  assign \U9_U2_U3_U0_DC_output[2] [14] = 1'b0;
  INV_X1_LVT U1_U0_U0_U1_i_0_0 (.A(A[4]), .ZN(\U1_U0_U0_U1_n_0[0] ));
  INV_X1_LVT U1_U0_U0_U1_i_0_1 (.A(B[19]), .ZN(\U1_U0_U0_U1_n_0[1] ));
  INV_X1_LVT U1_U0_U0_U1_i_0_2 (.A(U1_C[0]), .ZN(\U1_U0_U0_U1_n_0[2] ));
  OAI222_X1_LVT U1_U0_U0_U1_i_0_3 (.A1(\U1_U0_U0_U1_n_0[0] ), .A2(
      \U1_U0_U0_U1_n_0[1] ), .B1(\U1_U0_U0_U1_n_0[1] ), .B2(\U1_U0_U0_U1_n_0[2] ), 
      .C1(\U1_U0_U0_U1_n_0[0] ), .C2(\U1_U0_U0_U1_n_0[2] ), .ZN(U1_U0_C[1]));
  XNOR2_X1_LVT U1_U0_U0_U0_i_0_0 (.A(A[4]), .B(U1_C[0]), .ZN(
      \U1_U0_U0_U0_DC_output[1] [15]));
  XNOR2_X1_LVT U1_U0_U0_U0_i_0_1 (.A(\U1_U0_U0_U0_DC_output[1] [15]), .B(B[19]), 
      .ZN(SUM[2]));
  INV_X1_LVT U1_U0_U1_U1_i_0_0 (.A(A[5]), .ZN(\U1_U0_U1_U1_n_0[0] ));
  INV_X1_LVT U1_U0_U1_U1_i_0_1 (.A(B[20]), .ZN(\U1_U0_U1_U1_n_0[1] ));
  INV_X1_LVT U1_U0_U1_U1_i_0_2 (.A(U1_U0_C[1]), .ZN(\U1_U0_U1_U1_n_0[2] ));
  OAI222_X1_LVT U1_U0_U1_U1_i_0_3 (.A1(\U1_U0_U1_U1_n_0[0] ), .A2(
      \U1_U0_U1_U1_n_0[1] ), .B1(\U1_U0_U1_U1_n_0[1] ), .B2(\U1_U0_U1_U1_n_0[2] ), 
      .C1(\U1_U0_U1_U1_n_0[0] ), .C2(\U1_U0_U1_U1_n_0[2] ), .ZN(U1_U0_C[2]));
  XNOR2_X1_LVT U1_U0_U1_U0_i_0_0 (.A(A[5]), .B(U1_U0_C[1]), .ZN(
      \U1_U0_U1_U0_DC_output[1] [15]));
  XNOR2_X1_LVT U1_U0_U1_U0_i_0_1 (.A(\U1_U0_U1_U0_DC_output[1] [15]), .B(B[20]), 
      .ZN(SUM[3]));
  INV_X1_LVT U1_U0_U2_U1_i_0_0 (.A(A[6]), .ZN(\U1_U0_U2_U1_n_0[0] ));
  INV_X1_LVT U1_U0_U2_U1_i_0_1 (.A(B[21]), .ZN(\U1_U0_U2_U1_n_0[1] ));
  INV_X1_LVT U1_U0_U2_U1_i_0_2 (.A(U1_U0_C[2]), .ZN(\U1_U0_U2_U1_n_0[2] ));
  OAI222_X1_LVT U1_U0_U2_U1_i_0_3 (.A1(\U1_U0_U2_U1_n_0[0] ), .A2(
      \U1_U0_U2_U1_n_0[1] ), .B1(\U1_U0_U2_U1_n_0[1] ), .B2(\U1_U0_U2_U1_n_0[2] ), 
      .C1(\U1_U0_U2_U1_n_0[0] ), .C2(\U1_U0_U2_U1_n_0[2] ), .ZN(U1_U0_C[3]));
  XNOR2_X1_LVT U1_U0_U2_U0_i_0_0 (.A(A[6]), .B(U1_U0_C[2]), .ZN(
      \U1_U0_U2_U0_DC_output[1] [15]));
  XNOR2_X1_LVT U1_U0_U2_U0_i_0_1 (.A(\U1_U0_U2_U0_DC_output[1] [15]), .B(B[21]), 
      .ZN(SUM[4]));
  INV_X1_LVT U1_U0_U3_U1_i_0_0 (.A(A[7]), .ZN(\U1_U0_U3_U1_n_0[0] ));
  INV_X1_LVT U1_U0_U3_U1_i_0_1 (.A(B[22]), .ZN(\U1_U0_U3_U1_n_0[1] ));
  INV_X1_LVT U1_U0_U3_U1_i_0_2 (.A(U1_U0_C[3]), .ZN(\U1_U0_U3_U1_n_0[2] ));
  OAI222_X1_LVT U1_U0_U3_U1_i_0_3 (.A1(\U1_U0_U3_U1_n_0[0] ), .A2(
      \U1_U0_U3_U1_n_0[1] ), .B1(\U1_U0_U3_U1_n_0[1] ), .B2(\U1_U0_U3_U1_n_0[2] ), 
      .C1(\U1_U0_U3_U1_n_0[0] ), .C2(\U1_U0_U3_U1_n_0[2] ), .ZN(U1_C[1]));
  XNOR2_X1_LVT U1_U0_U3_U0_i_0_0 (.A(A[7]), .B(U1_U0_C[3]), .ZN(
      \U1_U0_U3_U0_DC_output[1] [15]));
  XNOR2_X1_LVT U1_U0_U3_U0_i_0_1 (.A(\U1_U0_U3_U0_DC_output[1] [15]), .B(B[22]), 
      .ZN(SUM[5]));
  INV_X1_LVT U1_U1_U0_U1_i_0_0 (.A(A[8]), .ZN(\U1_U1_U0_U1_n_0[0] ));
  INV_X1_LVT U1_U1_U0_U1_i_0_1 (.A(B[9]), .ZN(\U1_U1_U0_U1_n_0[1] ));
  INV_X1_LVT U1_U1_U0_U1_i_0_2 (.A(U1_C[1]), .ZN(\U1_U1_U0_U1_n_0[2] ));
  OAI222_X1_LVT U1_U1_U0_U1_i_0_3 (.A1(\U1_U1_U0_U1_n_0[0] ), .A2(
      \U1_U1_U0_U1_n_0[1] ), .B1(\U1_U1_U0_U1_n_0[1] ), .B2(\U1_U1_U0_U1_n_0[2] ), 
      .C1(\U1_U1_U0_U1_n_0[0] ), .C2(\U1_U1_U0_U1_n_0[2] ), .ZN(U1_U1_C[1]));
  XNOR2_X1_LVT U1_U1_U0_U0_i_0_0 (.A(A[8]), .B(U1_C[1]), .ZN(
      \U1_U1_U0_U0_DC_output[1] [15]));
  XNOR2_X1_LVT U1_U1_U0_U0_i_0_1 (.A(\U1_U1_U0_U0_DC_output[1] [15]), .B(B[9]), 
      .ZN(SUM[6]));
  INV_X1_LVT U1_U1_U1_U1_i_0_0 (.A(1'b0), .ZN(\U1_U1_U1_U1_n_0[0] ));
  INV_X1_LVT U1_U1_U1_U1_i_0_1 (.A(B[10]), .ZN(\U1_U1_U1_U1_n_0[1] ));
  INV_X1_LVT U1_U1_U1_U1_i_0_2 (.A(U1_U1_C[1]), .ZN(\U1_U1_U1_U1_n_0[2] ));
  OAI222_X1_LVT U1_U1_U1_U1_i_0_3 (.A1(\U1_U1_U1_U1_n_0[0] ), .A2(
      \U1_U1_U1_U1_n_0[1] ), .B1(\U1_U1_U1_U1_n_0[1] ), .B2(\U1_U1_U1_U1_n_0[2] ), 
      .C1(\U1_U1_U1_U1_n_0[0] ), .C2(\U1_U1_U1_U1_n_0[2] ), .ZN(U1_U1_C[2]));
  XNOR2_X1_LVT U1_U1_U1_U0_i_0_0 (.A(1'b0), .B(U1_U1_C[1]), .ZN(
      \U1_U1_U1_U0_DC_output[1] [15]));
  XNOR2_X1_LVT U1_U1_U1_U0_i_0_1 (.A(\U1_U1_U1_U0_DC_output[1] [15]), .B(B[10]), 
      .ZN(SUM[7]));
  INV_X1_LVT U1_U1_U2_U1_i_0_0 (.A(A[3]), .ZN(\U1_U1_U2_U1_n_0[0] ));
  INV_X1_LVT U1_U1_U2_U1_i_0_1 (.A(B[11]), .ZN(\U1_U1_U2_U1_n_0[1] ));
  INV_X1_LVT U1_U1_U2_U1_i_0_2 (.A(U1_U1_C[2]), .ZN(\U1_U1_U2_U1_n_0[2] ));
  OAI222_X1_LVT U1_U1_U2_U1_i_0_3 (.A1(\U1_U1_U2_U1_n_0[0] ), .A2(
      \U1_U1_U2_U1_n_0[1] ), .B1(\U1_U1_U2_U1_n_0[1] ), .B2(\U1_U1_U2_U1_n_0[2] ), 
      .C1(\U1_U1_U2_U1_n_0[0] ), .C2(\U1_U1_U2_U1_n_0[2] ), .ZN(U1_U1_C[3]));
  XNOR2_X1_LVT U1_U1_U2_U0_i_0_0 (.A(A[3]), .B(U1_U1_C[2]), .ZN(
      \U1_U1_U2_U0_DC_output[1] [15]));
  XNOR2_X1_LVT U1_U1_U2_U0_i_0_1 (.A(\U1_U1_U2_U0_DC_output[1] [15]), .B(B[11]), 
      .ZN(SUM[8]));
  INV_X1_LVT U1_U1_U3_U1_i_0_0 (.A(A[1]), .ZN(\U1_U1_U3_U1_n_0[0] ));
  INV_X1_LVT U1_U1_U3_U1_i_0_1 (.A(B[0]), .ZN(\U1_U1_U3_U1_n_0[1] ));
  INV_X1_LVT U1_U1_U3_U1_i_0_2 (.A(U1_U1_C[3]), .ZN(\U1_U1_U3_U1_n_0[2] ));
  OAI222_X1_LVT U1_U1_U3_U1_i_0_3 (.A1(\U1_U1_U3_U1_n_0[0] ), .A2(
      \U1_U1_U3_U1_n_0[1] ), .B1(\U1_U1_U3_U1_n_0[1] ), .B2(\U1_U1_U3_U1_n_0[2] ), 
      .C1(\U1_U1_U3_U1_n_0[0] ), .C2(\U1_U1_U3_U1_n_0[2] ), .ZN(U1_C[2]));
  XNOR2_X1_LVT U1_U1_U3_U0_i_0_0 (.A(A[1]), .B(U1_U1_C[3]), .ZN(
      \U1_U1_U3_U0_DC_output[1] [15]));
  XNOR2_X1_LVT U1_U1_U3_U0_i_0_1 (.A(\U1_U1_U3_U0_DC_output[1] [15]), .B(B[0]), 
      .ZN(SUM[9]));
  INV_X1_LVT U1_U2_U0_U1_i_0_0 (.A(1'b1), .ZN(\U1_U2_U0_U1_n_0[0] ));
  INV_X1_LVT U1_U2_U0_U1_i_0_1 (.A(1'b1), .ZN(\U1_U2_U0_U1_n_0[1] ));
  INV_X1_LVT U1_U2_U0_U1_i_0_2 (.A(U1_C[2]), .ZN(\U1_U2_U0_U1_n_0[2] ));
  OAI222_X1_LVT U1_U2_U0_U1_i_0_3 (.A1(\U1_U2_U0_U1_n_0[0] ), .A2(
      \U1_U2_U0_U1_n_0[1] ), .B1(\U1_U2_U0_U1_n_0[1] ), .B2(\U1_U2_U0_U1_n_0[2] ), 
      .C1(\U1_U2_U0_U1_n_0[0] ), .C2(\U1_U2_U0_U1_n_0[2] ), .ZN(U1_U2_C[1]));
  XNOR2_X1_LVT U1_U2_U0_U0_i_0_0 (.A(1'b1), .B(U1_C[2]), .ZN(
      \U1_U2_U0_U0_DC_output[1] [15]));
  XNOR2_X1_LVT U1_U2_U0_U0_i_0_1 (.A(\U1_U2_U0_U0_DC_output[1] [15]), .B(1'b1), 
      .ZN(SUM[10]));
  INV_X1_LVT U1_U2_U1_U1_i_0_0 (.A(1'b0), .ZN(\U1_U2_U1_U1_n_0[0] ));
  INV_X1_LVT U1_U2_U1_U1_i_0_1 (.A(1'b1), .ZN(\U1_U2_U1_U1_n_0[1] ));
  INV_X1_LVT U1_U2_U1_U1_i_0_2 (.A(U1_U2_C[1]), .ZN(\U1_U2_U1_U1_n_0[2] ));
  OAI222_X1_LVT U1_U2_U1_U1_i_0_3 (.A1(\U1_U2_U1_U1_n_0[0] ), .A2(
      \U1_U2_U1_U1_n_0[1] ), .B1(\U1_U2_U1_U1_n_0[1] ), .B2(\U1_U2_U1_U1_n_0[2] ), 
      .C1(\U1_U2_U1_U1_n_0[0] ), .C2(\U1_U2_U1_U1_n_0[2] ), .ZN(U1_U2_C[2]));
  XNOR2_X1_LVT U1_U2_U1_U0_i_0_0 (.A(1'b0), .B(U1_U2_C[1]), .ZN(
      \U1_U2_U1_U0_DC_output[1] [15]));
  XNOR2_X1_LVT U1_U2_U1_U0_i_0_1 (.A(\U1_U2_U1_U0_DC_output[1] [15]), .B(1'b1), 
      .ZN(SUM[11]));
  INV_X1_LVT U1_U2_U2_U1_i_0_0 (.A(1'b1), .ZN(\U1_U2_U2_U1_n_0[0] ));
  INV_X1_LVT U1_U2_U2_U1_i_0_1 (.A(1'b0), .ZN(\U1_U2_U2_U1_n_0[1] ));
  INV_X1_LVT U1_U2_U2_U1_i_0_2 (.A(U1_U2_C[2]), .ZN(\U1_U2_U2_U1_n_0[2] ));
  OAI222_X1_LVT U1_U2_U2_U1_i_0_3 (.A1(\U1_U2_U2_U1_n_0[0] ), .A2(
      \U1_U2_U2_U1_n_0[1] ), .B1(\U1_U2_U2_U1_n_0[1] ), .B2(\U1_U2_U2_U1_n_0[2] ), 
      .C1(\U1_U2_U2_U1_n_0[0] ), .C2(\U1_U2_U2_U1_n_0[2] ), .ZN(U1_U2_C[3]));
  XNOR2_X1_LVT U1_U2_U2_U0_i_0_0 (.A(1'b1), .B(U1_U2_C[2]), .ZN(
      \U1_U2_U2_U0_DC_output[1] [15]));
  XNOR2_X1_LVT U1_U2_U2_U0_i_0_1 (.A(\U1_U2_U2_U0_DC_output[1] [15]), .B(1'b0), 
      .ZN(SUM[12]));
  INV_X1_LVT U1_U2_U3_U1_i_0_0 (.A(1'b0), .ZN(\U1_U2_U3_U1_n_0[0] ));
  INV_X1_LVT U1_U2_U3_U1_i_0_1 (.A(1'b0), .ZN(\U1_U2_U3_U1_n_0[1] ));
  INV_X1_LVT U1_U2_U3_U1_i_0_2 (.A(U1_U2_C[3]), .ZN(\U1_U2_U3_U1_n_0[2] ));
  OAI222_X1_LVT U1_U2_U3_U1_i_0_3 (.A1(\U1_U2_U3_U1_n_0[0] ), .A2(
      \U1_U2_U3_U1_n_0[1] ), .B1(\U1_U2_U3_U1_n_0[1] ), .B2(\U1_U2_U3_U1_n_0[2] ), 
      .C1(\U1_U2_U3_U1_n_0[0] ), .C2(\U1_U2_U3_U1_n_0[2] ), .ZN(U1_c_no_defined));
  XNOR2_X1_LVT U1_U2_U3_U0_i_0_0 (.A(1'b0), .B(U1_U2_C[3]), .ZN(
      \U1_U2_U3_U0_DC_output[1] [15]));
  XNOR2_X1_LVT U1_U2_U3_U0_i_0_1 (.A(\U1_U2_U3_U0_DC_output[1] [15]), .B(1'b0), 
      .ZN(SUM[13]));
  INV_X1_LVT U2_U0_U0_U1_i_0_0 (.A(A[9]), .ZN(\U2_U0_U0_U1_n_0[0] ));
  INV_X1_LVT U2_U0_U0_U1_i_0_1 (.A(B[12]), .ZN(\U2_U0_U0_U1_n_0[1] ));
  INV_X1_LVT U2_U0_U0_U1_i_0_2 (.A(U2_C[0]), .ZN(\U2_U0_U0_U1_n_0[2] ));
  OAI222_X1_LVT U2_U0_U0_U1_i_0_3 (.A1(\U2_U0_U0_U1_n_0[0] ), .A2(
      \U2_U0_U0_U1_n_0[1] ), .B1(\U2_U0_U0_U1_n_0[1] ), .B2(\U2_U0_U0_U1_n_0[2] ), 
      .C1(\U2_U0_U0_U1_n_0[0] ), .C2(\U2_U0_U0_U1_n_0[2] ), .ZN(U2_U0_C[1]));
  XNOR2_X1_LVT U2_U0_U0_U0_i_0_0 (.A(A[9]), .B(U2_C[0]), .ZN(
      \U2_U0_U0_U0_DC_output[1] [15]));
  XNOR2_X1_LVT U2_U0_U0_U0_i_0_1 (.A(\U2_U0_U0_U0_DC_output[1] [15]), .B(B[12]), 
      .ZN(SUM[14]));
  INV_X1_LVT U2_U0_U1_U1_i_0_0 (.A(A[10]), .ZN(\U2_U0_U1_U1_n_0[0] ));
  INV_X1_LVT U2_U0_U1_U1_i_0_1 (.A(B[13]), .ZN(\U2_U0_U1_U1_n_0[1] ));
  INV_X1_LVT U2_U0_U1_U1_i_0_2 (.A(U2_U0_C[1]), .ZN(\U2_U0_U1_U1_n_0[2] ));
  OAI222_X1_LVT U2_U0_U1_U1_i_0_3 (.A1(\U2_U0_U1_U1_n_0[0] ), .A2(
      \U2_U0_U1_U1_n_0[1] ), .B1(\U2_U0_U1_U1_n_0[1] ), .B2(\U2_U0_U1_U1_n_0[2] ), 
      .C1(\U2_U0_U1_U1_n_0[0] ), .C2(\U2_U0_U1_U1_n_0[2] ), .ZN(U2_U0_C[2]));
  XNOR2_X1_LVT U2_U0_U1_U0_i_0_0 (.A(A[10]), .B(U2_U0_C[1]), .ZN(
      \U2_U0_U1_U0_DC_output[1] [15]));
  XNOR2_X1_LVT U2_U0_U1_U0_i_0_1 (.A(\U2_U0_U1_U0_DC_output[1] [15]), .B(B[13]), 
      .ZN(SUM[15]));
  INV_X1_LVT U2_U0_U2_U1_i_0_0 (.A(A[11]), .ZN(\U2_U0_U2_U1_n_0[0] ));
  INV_X1_LVT U2_U0_U2_U1_i_0_1 (.A(B[14]), .ZN(\U2_U0_U2_U1_n_0[1] ));
  INV_X1_LVT U2_U0_U2_U1_i_0_2 (.A(U2_U0_C[2]), .ZN(\U2_U0_U2_U1_n_0[2] ));
  OAI222_X1_LVT U2_U0_U2_U1_i_0_3 (.A1(\U2_U0_U2_U1_n_0[0] ), .A2(
      \U2_U0_U2_U1_n_0[1] ), .B1(\U2_U0_U2_U1_n_0[1] ), .B2(\U2_U0_U2_U1_n_0[2] ), 
      .C1(\U2_U0_U2_U1_n_0[0] ), .C2(\U2_U0_U2_U1_n_0[2] ), .ZN(U2_U0_C[3]));
  XNOR2_X1_LVT U2_U0_U2_U0_i_0_0 (.A(A[11]), .B(U2_U0_C[2]), .ZN(
      \U2_U0_U2_U0_DC_output[1] [15]));
  XNOR2_X1_LVT U2_U0_U2_U0_i_0_1 (.A(\U2_U0_U2_U0_DC_output[1] [15]), .B(B[14]), 
      .ZN(SUM[16]));
  INV_X1_LVT U2_U0_U3_U1_i_0_0 (.A(A[12]), .ZN(\U2_U0_U3_U1_n_0[0] ));
  INV_X1_LVT U2_U0_U3_U1_i_0_1 (.A(B[15]), .ZN(\U2_U0_U3_U1_n_0[1] ));
  INV_X1_LVT U2_U0_U3_U1_i_0_2 (.A(U2_U0_C[3]), .ZN(\U2_U0_U3_U1_n_0[2] ));
  OAI222_X1_LVT U2_U0_U3_U1_i_0_3 (.A1(\U2_U0_U3_U1_n_0[0] ), .A2(
      \U2_U0_U3_U1_n_0[1] ), .B1(\U2_U0_U3_U1_n_0[1] ), .B2(\U2_U0_U3_U1_n_0[2] ), 
      .C1(\U2_U0_U3_U1_n_0[0] ), .C2(\U2_U0_U3_U1_n_0[2] ), .ZN(U2_C[1]));
  XNOR2_X1_LVT U2_U0_U3_U0_i_0_0 (.A(A[12]), .B(U2_U0_C[3]), .ZN(
      \U2_U0_U3_U0_DC_output[1] [15]));
  XNOR2_X1_LVT U2_U0_U3_U0_i_0_1 (.A(\U2_U0_U3_U0_DC_output[1] [15]), .B(B[15]), 
      .ZN(SUM[17]));
  INV_X1_LVT U2_U1_U0_U1_i_0_0 (.A(A[13]), .ZN(\U2_U1_U0_U1_n_0[0] ));
  INV_X1_LVT U2_U1_U0_U1_i_0_1 (.A(B[16]), .ZN(\U2_U1_U0_U1_n_0[1] ));
  INV_X1_LVT U2_U1_U0_U1_i_0_2 (.A(U2_C[1]), .ZN(\U2_U1_U0_U1_n_0[2] ));
  OAI222_X1_LVT U2_U1_U0_U1_i_0_3 (.A1(\U2_U1_U0_U1_n_0[0] ), .A2(
      \U2_U1_U0_U1_n_0[1] ), .B1(\U2_U1_U0_U1_n_0[1] ), .B2(\U2_U1_U0_U1_n_0[2] ), 
      .C1(\U2_U1_U0_U1_n_0[0] ), .C2(\U2_U1_U0_U1_n_0[2] ), .ZN(U2_U1_C[1]));
  XNOR2_X1_LVT U2_U1_U0_U0_i_0_0 (.A(A[13]), .B(U2_C[1]), .ZN(
      \U2_U1_U0_U0_DC_output[1] [15]));
  XNOR2_X1_LVT U2_U1_U0_U0_i_0_1 (.A(\U2_U1_U0_U0_DC_output[1] [15]), .B(B[16]), 
      .ZN(SUM[18]));
  INV_X1_LVT U2_U1_U1_U1_i_0_0 (.A(A[14]), .ZN(\U2_U1_U1_U1_n_0[0] ));
  INV_X1_LVT U2_U1_U1_U1_i_0_1 (.A(B[17]), .ZN(\U2_U1_U1_U1_n_0[1] ));
  INV_X1_LVT U2_U1_U1_U1_i_0_2 (.A(U2_U1_C[1]), .ZN(\U2_U1_U1_U1_n_0[2] ));
  OAI222_X1_LVT U2_U1_U1_U1_i_0_3 (.A1(\U2_U1_U1_U1_n_0[0] ), .A2(
      \U2_U1_U1_U1_n_0[1] ), .B1(\U2_U1_U1_U1_n_0[1] ), .B2(\U2_U1_U1_U1_n_0[2] ), 
      .C1(\U2_U1_U1_U1_n_0[0] ), .C2(\U2_U1_U1_U1_n_0[2] ), .ZN(U2_U1_C[2]));
  XNOR2_X1_LVT U2_U1_U1_U0_i_0_0 (.A(A[14]), .B(U2_U1_C[1]), .ZN(
      \U2_U1_U1_U0_DC_output[1] [15]));
  XNOR2_X1_LVT U2_U1_U1_U0_i_0_1 (.A(\U2_U1_U1_U0_DC_output[1] [15]), .B(B[17]), 
      .ZN(SUM[19]));
  INV_X1_LVT U2_U1_U2_U1_i_0_0 (.A(A[15]), .ZN(\U2_U1_U2_U1_n_0[0] ));
  INV_X1_LVT U2_U1_U2_U1_i_0_1 (.A(B[18]), .ZN(\U2_U1_U2_U1_n_0[1] ));
  INV_X1_LVT U2_U1_U2_U1_i_0_2 (.A(U2_U1_C[2]), .ZN(\U2_U1_U2_U1_n_0[2] ));
  OAI222_X1_LVT U2_U1_U2_U1_i_0_3 (.A1(\U2_U1_U2_U1_n_0[0] ), .A2(
      \U2_U1_U2_U1_n_0[1] ), .B1(\U2_U1_U2_U1_n_0[1] ), .B2(\U2_U1_U2_U1_n_0[2] ), 
      .C1(\U2_U1_U2_U1_n_0[0] ), .C2(\U2_U1_U2_U1_n_0[2] ), .ZN(U2_U1_C[3]));
  XNOR2_X1_LVT U2_U1_U2_U0_i_0_0 (.A(A[15]), .B(U2_U1_C[2]), .ZN(
      \U2_U1_U2_U0_DC_output[1] [15]));
  XNOR2_X1_LVT U2_U1_U2_U0_i_0_1 (.A(\U2_U1_U2_U0_DC_output[1] [15]), .B(B[18]), 
      .ZN(SUM[20]));
  INV_X1_LVT U2_U1_U3_U1_i_0_0 (.A(A[16]), .ZN(\U2_U1_U3_U1_n_0[0] ));
  INV_X1_LVT U2_U1_U3_U1_i_0_1 (.A(B[4]), .ZN(\U2_U1_U3_U1_n_0[1] ));
  INV_X1_LVT U2_U1_U3_U1_i_0_2 (.A(U2_U1_C[3]), .ZN(\U2_U1_U3_U1_n_0[2] ));
  OAI222_X1_LVT U2_U1_U3_U1_i_0_3 (.A1(\U2_U1_U3_U1_n_0[0] ), .A2(
      \U2_U1_U3_U1_n_0[1] ), .B1(\U2_U1_U3_U1_n_0[1] ), .B2(\U2_U1_U3_U1_n_0[2] ), 
      .C1(\U2_U1_U3_U1_n_0[0] ), .C2(\U2_U1_U3_U1_n_0[2] ), .ZN(U2_C[2]));
  XNOR2_X1_LVT U2_U1_U3_U0_i_0_0 (.A(A[16]), .B(U2_U1_C[3]), .ZN(
      \U2_U1_U3_U0_DC_output[1] [15]));
  XNOR2_X1_LVT U2_U1_U3_U0_i_0_1 (.A(\U2_U1_U3_U0_DC_output[1] [15]), .B(B[4]), 
      .ZN(SUM[21]));
  INV_X1_LVT U2_U2_U0_U1_i_0_0 (.A(A[17]), .ZN(\U2_U2_U0_U1_n_0[0] ));
  INV_X1_LVT U2_U2_U0_U1_i_0_1 (.A(B[5]), .ZN(\U2_U2_U0_U1_n_0[1] ));
  INV_X1_LVT U2_U2_U0_U1_i_0_2 (.A(U2_C[2]), .ZN(\U2_U2_U0_U1_n_0[2] ));
  OAI222_X1_LVT U2_U2_U0_U1_i_0_3 (.A1(\U2_U2_U0_U1_n_0[0] ), .A2(
      \U2_U2_U0_U1_n_0[1] ), .B1(\U2_U2_U0_U1_n_0[1] ), .B2(\U2_U2_U0_U1_n_0[2] ), 
      .C1(\U2_U2_U0_U1_n_0[0] ), .C2(\U2_U2_U0_U1_n_0[2] ), .ZN(U2_U2_C[1]));
  XNOR2_X1_LVT U2_U2_U0_U0_i_0_0 (.A(A[17]), .B(U2_C[2]), .ZN(
      \U2_U2_U0_U0_DC_output[1] [15]));
  XNOR2_X1_LVT U2_U2_U0_U0_i_0_1 (.A(\U2_U2_U0_U0_DC_output[1] [15]), .B(B[5]), 
      .ZN(SUM[22]));
  INV_X1_LVT U2_U2_U1_U1_i_0_0 (.A(A[18]), .ZN(\U2_U2_U1_U1_n_0[0] ));
  INV_X1_LVT U2_U2_U1_U1_i_0_1 (.A(B[6]), .ZN(\U2_U2_U1_U1_n_0[1] ));
  INV_X1_LVT U2_U2_U1_U1_i_0_2 (.A(U2_U2_C[1]), .ZN(\U2_U2_U1_U1_n_0[2] ));
  OAI222_X1_LVT U2_U2_U1_U1_i_0_3 (.A1(\U2_U2_U1_U1_n_0[0] ), .A2(
      \U2_U2_U1_U1_n_0[1] ), .B1(\U2_U2_U1_U1_n_0[1] ), .B2(\U2_U2_U1_U1_n_0[2] ), 
      .C1(\U2_U2_U1_U1_n_0[0] ), .C2(\U2_U2_U1_U1_n_0[2] ), .ZN(U2_U2_C[2]));
  XNOR2_X1_LVT U2_U2_U1_U0_i_0_0 (.A(A[18]), .B(U2_U2_C[1]), .ZN(
      \U2_U2_U1_U0_DC_output[1] [15]));
  XNOR2_X1_LVT U2_U2_U1_U0_i_0_1 (.A(\U2_U2_U1_U0_DC_output[1] [15]), .B(B[6]), 
      .ZN(SUM[23]));
  INV_X1_LVT U2_U2_U2_U1_i_0_0 (.A(A[2]), .ZN(\U2_U2_U2_U1_n_0[0] ));
  INV_X1_LVT U2_U2_U2_U1_i_0_1 (.A(B[7]), .ZN(\U2_U2_U2_U1_n_0[1] ));
  INV_X1_LVT U2_U2_U2_U1_i_0_2 (.A(U2_U2_C[2]), .ZN(\U2_U2_U2_U1_n_0[2] ));
  OAI222_X1_LVT U2_U2_U2_U1_i_0_3 (.A1(\U2_U2_U2_U1_n_0[0] ), .A2(
      \U2_U2_U2_U1_n_0[1] ), .B1(\U2_U2_U2_U1_n_0[1] ), .B2(\U2_U2_U2_U1_n_0[2] ), 
      .C1(\U2_U2_U2_U1_n_0[0] ), .C2(\U2_U2_U2_U1_n_0[2] ), .ZN(U2_U2_C[3]));
  XNOR2_X1_LVT U2_U2_U2_U0_i_0_0 (.A(A[2]), .B(U2_U2_C[2]), .ZN(
      \U2_U2_U2_U0_DC_output[1] [15]));
  XNOR2_X1_LVT U2_U2_U2_U0_i_0_1 (.A(\U2_U2_U2_U0_DC_output[1] [15]), .B(B[7]), 
      .ZN(SUM[24]));
  INV_X1_LVT U2_U2_U3_U1_i_0_0 (.A(A[0]), .ZN(\U2_U2_U3_U1_n_0[0] ));
  INV_X1_LVT U2_U2_U3_U1_i_0_1 (.A(B[8]), .ZN(\U2_U2_U3_U1_n_0[1] ));
  INV_X1_LVT U2_U2_U3_U1_i_0_2 (.A(U2_U2_C[3]), .ZN(\U2_U2_U3_U1_n_0[2] ));
  OAI222_X1_LVT U2_U2_U3_U1_i_0_3 (.A1(\U2_U2_U3_U1_n_0[0] ), .A2(
      \U2_U2_U3_U1_n_0[1] ), .B1(\U2_U2_U3_U1_n_0[1] ), .B2(\U2_U2_U3_U1_n_0[2] ), 
      .C1(\U2_U2_U3_U1_n_0[0] ), .C2(\U2_U2_U3_U1_n_0[2] ), .ZN(U2_c_no_defined));
  XNOR2_X1_LVT U2_U2_U3_U0_i_0_0 (.A(A[0]), .B(U2_U2_C[3]), .ZN(
      \U2_U2_U3_U0_DC_output[1] [15]));
  XNOR2_X1_LVT U2_U2_U3_U0_i_0_1 (.A(\U2_U2_U3_U0_DC_output[1] [15]), .B(B[8]), 
      .ZN(SUM[25]));
  INV_X1_LVT U3_U1_i_0_0 (.A(1'b1), .ZN(\U3_U1_n_0[0] ));
  INV_X1_LVT U3_U1_i_0_1 (.A(1'b0), .ZN(\U3_U1_n_0[1] ));
  INV_X1_LVT U3_U1_i_0_2 (.A(C[2]), .ZN(\U3_U1_n_0[2] ));
  OAI222_X1_LVT U3_U1_i_0_3 (.A1(\U3_U1_n_0[0] ), .A2(\U3_U1_n_0[1] ), .B1(
      \U3_U1_n_0[1] ), .B2(\U3_U1_n_0[2] ), .C1(\U3_U1_n_0[0] ), .C2(
      \U3_U1_n_0[2] ), .ZN(C[1]));
  XNOR2_X1_LVT U3_U0_i_0_0 (.A(1'b1), .B(C[2]), .ZN(\U3_U0_DC_output[1] [15]));
  XNOR2_X1_LVT U3_U0_i_0_1 (.A(\U3_U0_DC_output[1] [15]), .B(1'b0), .ZN(SUM[0]));
  INV_X1_LVT U4_U1_i_0_0 (.A(C[0]), .ZN(\U4_U1_n_0[0] ));
  INV_X1_LVT U4_U1_i_0_1 (.A(C[3]), .ZN(\U4_U1_n_0[1] ));
  INV_X1_LVT U4_U1_i_0_2 (.A(C[1]), .ZN(\U4_U1_n_0[2] ));
  OAI222_X1_LVT U4_U1_i_0_3 (.A1(\U4_U1_n_0[0] ), .A2(\U4_U1_n_0[1] ), .B1(
      \U4_U1_n_0[1] ), .B2(\U4_U1_n_0[2] ), .C1(\U4_U1_n_0[0] ), .C2(
      \U4_U1_n_0[2] ), .ZN(C[9]));
  XNOR2_X1_LVT U4_U0_i_0_0 (.A(C[0]), .B(C[1]), .ZN(\U4_U0_DC_output[1] [15]));
  XNOR2_X1_LVT U4_U0_i_0_1 (.A(\U4_U0_DC_output[1] [15]), .B(C[3]), .ZN(SUM[1]));
  INV_X1_LVT U5_i_0_0 (.A(A[23]), .ZN(\U5_n_0[0] ));
  INV_X1_LVT U5_i_0_1 (.A(B[23]), .ZN(\U5_n_0[1] ));
  INV_X1_LVT U5_i_0_2 (.A(cci), .ZN(\U5_n_0[2] ));
  OAI222_X1_LVT U5_i_0_3 (.A1(\U5_n_0[0] ), .A2(\U5_n_0[1] ), .B1(\U5_n_0[1] ), 
      .B2(\U5_n_0[2] ), .C1(\U5_n_0[0] ), .C2(\U5_n_0[2] ), .ZN(C[7]));
  INV_X1_LVT U6_U0_U1_i_0_0 (.A(A[19]), .ZN(\U6_U0_U1_n_0[0] ));
  INV_X1_LVT U6_U0_U1_i_0_1 (.A(1'b1), .ZN(\U6_U0_U1_n_0[1] ));
  INV_X1_LVT U6_U0_U1_i_0_2 (.A(C[0]), .ZN(\U6_U0_U1_n_0[2] ));
  OAI222_X1_LVT U6_U0_U1_i_0_3 (.A1(\U6_U0_U1_n_0[0] ), .A2(\U6_U0_U1_n_0[1] ), 
      .B1(\U6_U0_U1_n_0[1] ), .B2(\U6_U0_U1_n_0[2] ), .C1(\U6_U0_U1_n_0[0] ), 
      .C2(\U6_U0_U1_n_0[2] ), .ZN(U6_C[1]));
  XNOR2_X1_LVT U6_U0_U0_i_0_0 (.A(A[19]), .B(C[0]), .ZN(\U6_U0_U0_DC_output[1] [15]));
  XNOR2_X1_LVT U6_U0_U0_i_0_1 (.A(\U6_U0_U0_DC_output[1] [15]), .B(1'b1), .ZN(
      SUM[26]));
  INV_X1_LVT U6_U1_U1_i_0_0 (.A(A[20]), .ZN(\U6_U1_U1_n_0[0] ));
  INV_X1_LVT U6_U1_U1_i_0_1 (.A(B[1]), .ZN(\U6_U1_U1_n_0[1] ));
  INV_X1_LVT U6_U1_U1_i_0_2 (.A(U6_C[1]), .ZN(\U6_U1_U1_n_0[2] ));
  OAI222_X1_LVT U6_U1_U1_i_0_3 (.A1(\U6_U1_U1_n_0[0] ), .A2(\U6_U1_U1_n_0[1] ), 
      .B1(\U6_U1_U1_n_0[1] ), .B2(\U6_U1_U1_n_0[2] ), .C1(\U6_U1_U1_n_0[0] ), 
      .C2(\U6_U1_U1_n_0[2] ), .ZN(U6_C[2]));
  XNOR2_X1_LVT U6_U1_U0_i_0_0 (.A(A[20]), .B(U6_C[1]), .ZN(
      \U6_U1_U0_DC_output[1] [15]));
  XNOR2_X1_LVT U6_U1_U0_i_0_1 (.A(\U6_U1_U0_DC_output[1] [15]), .B(B[1]), .ZN(
      SUM[27]));
  INV_X1_LVT U6_U2_U1_i_0_0 (.A(A[21]), .ZN(\U6_U2_U1_n_0[0] ));
  INV_X1_LVT U6_U2_U1_i_0_1 (.A(B[2]), .ZN(\U6_U2_U1_n_0[1] ));
  INV_X1_LVT U6_U2_U1_i_0_2 (.A(U6_C[2]), .ZN(\U6_U2_U1_n_0[2] ));
  OAI222_X1_LVT U6_U2_U1_i_0_3 (.A1(\U6_U2_U1_n_0[0] ), .A2(\U6_U2_U1_n_0[1] ), 
      .B1(\U6_U2_U1_n_0[1] ), .B2(\U6_U2_U1_n_0[2] ), .C1(\U6_U2_U1_n_0[0] ), 
      .C2(\U6_U2_U1_n_0[2] ), .ZN(U6_C[3]));
  XNOR2_X1_LVT U6_U2_U0_i_0_0 (.A(A[21]), .B(U6_C[2]), .ZN(
      \U6_U2_U0_DC_output[1] [15]));
  XNOR2_X1_LVT U6_U2_U0_i_0_1 (.A(\U6_U2_U0_DC_output[1] [15]), .B(B[2]), .ZN(
      SUM[28]));
  INV_X1_LVT U6_U3_U1_i_0_0 (.A(A[22]), .ZN(\U6_U3_U1_n_0[0] ));
  INV_X1_LVT U6_U3_U1_i_0_1 (.A(B[3]), .ZN(\U6_U3_U1_n_0[1] ));
  INV_X1_LVT U6_U3_U1_i_0_2 (.A(U6_C[3]), .ZN(\U6_U3_U1_n_0[2] ));
  OAI222_X1_LVT U6_U3_U1_i_0_3 (.A1(\U6_U3_U1_n_0[0] ), .A2(\U6_U3_U1_n_0[1] ), 
      .B1(\U6_U3_U1_n_0[1] ), .B2(\U6_U3_U1_n_0[2] ), .C1(\U6_U3_U1_n_0[0] ), 
      .C2(\U6_U3_U1_n_0[2] ), .ZN(C[8]));
  XNOR2_X1_LVT U6_U3_U0_i_0_0 (.A(A[22]), .B(U6_C[3]), .ZN(
      \U6_U3_U0_DC_output[1] [15]));
  XNOR2_X1_LVT U6_U3_U0_i_0_1 (.A(\U6_U3_U0_DC_output[1] [15]), .B(B[3]), .ZN(
      SUM[29]));
  SDFF_X1_LVT U7 (.CK(1'b1), .D(), .SE(1'b0), .SI(1'b1), .Q(), .QN());
  INV_X1_LVT U8_U0_U1_i_0_0 (.A(1'b0), .ZN(\U8_U0_U1_n_0[0] ));
  INV_X1_LVT U8_U0_U1_i_0_1 (.A(1'b1), .ZN(\U8_U0_U1_n_0[1] ));
  INV_X1_LVT U8_U0_U1_i_0_2 (.A(), .ZN(\U8_U0_U1_n_0[2] ));
  OAI222_X1_LVT U8_U0_U1_i_0_3 (.A1(\U8_U0_U1_n_0[0] ), .A2(\U8_U0_U1_n_0[1] ), 
      .B1(\U8_U0_U1_n_0[1] ), .B2(\U8_U0_U1_n_0[2] ), .C1(\U8_U0_U1_n_0[0] ), 
      .C2(\U8_U0_U1_n_0[2] ), .ZN(U8_C[1]));
  XNOR2_X1_LVT U8_U0_U0_i_0_0 (.A(1'b0), .B(), .ZN(\U8_U0_U0_DC_output[1] [15]));
  XNOR2_X1_LVT U8_U0_U0_i_0_1 (.A(\U8_U0_U0_DC_output[1] [15]), .B(1'b1), .ZN());
  INV_X1_LVT U8_U1_U1_i_0_0 (.A(ci), .ZN(\U8_U1_U1_n_0[0] ));
  INV_X1_LVT U8_U1_U1_i_0_1 (.A(1'b1), .ZN(\U8_U1_U1_n_0[1] ));
  INV_X1_LVT U8_U1_U1_i_0_2 (.A(U8_C[1]), .ZN(\U8_U1_U1_n_0[2] ));
  OAI222_X1_LVT U8_U1_U1_i_0_3 (.A1(\U8_U1_U1_n_0[0] ), .A2(\U8_U1_U1_n_0[1] ), 
      .B1(\U8_U1_U1_n_0[1] ), .B2(\U8_U1_U1_n_0[2] ), .C1(\U8_U1_U1_n_0[0] ), 
      .C2(\U8_U1_U1_n_0[2] ), .ZN(U8_C[2]));
  XNOR2_X1_LVT U8_U1_U0_i_0_0 (.A(ci), .B(U8_C[1]), .ZN(
      \U8_U1_U0_DC_output[1] [15]));
  XNOR2_X1_LVT U8_U1_U0_i_0_1 (.A(\U8_U1_U0_DC_output[1] [15]), .B(1'b1), .ZN());
  INV_X1_LVT U8_U2_U1_i_0_0 (.A(1'b0), .ZN(\U8_U2_U1_n_0[0] ));
  INV_X1_LVT U8_U2_U1_i_0_1 (.A(ci), .ZN(\U8_U2_U1_n_0[1] ));
  INV_X1_LVT U8_U2_U1_i_0_2 (.A(U8_C[2]), .ZN(\U8_U2_U1_n_0[2] ));
  OAI222_X1_LVT U8_U2_U1_i_0_3 (.A1(\U8_U2_U1_n_0[0] ), .A2(\U8_U2_U1_n_0[1] ), 
      .B1(\U8_U2_U1_n_0[1] ), .B2(\U8_U2_U1_n_0[2] ), .C1(\U8_U2_U1_n_0[0] ), 
      .C2(\U8_U2_U1_n_0[2] ), .ZN(U8_C[3]));
  XNOR2_X1_LVT U8_U2_U0_i_0_0 (.A(1'b0), .B(U8_C[2]), .ZN(
      \U8_U2_U0_DC_output[1] [15]));
  XNOR2_X1_LVT U8_U2_U0_i_0_1 (.A(\U8_U2_U0_DC_output[1] [15]), .B(ci), .ZN());
  INV_X1_LVT U8_U3_U1_i_0_0 (.A(1'b0), .ZN(\U8_U3_U1_n_0[0] ));
  INV_X1_LVT U8_U3_U1_i_0_1 (.A(1'b0), .ZN(\U8_U3_U1_n_0[1] ));
  INV_X1_LVT U8_U3_U1_i_0_2 (.A(U8_C[3]), .ZN(\U8_U3_U1_n_0[2] ));
  OAI222_X1_LVT U8_U3_U1_i_0_3 (.A1(\U8_U3_U1_n_0[0] ), .A2(\U8_U3_U1_n_0[1] ), 
      .B1(\U8_U3_U1_n_0[1] ), .B2(\U8_U3_U1_n_0[2] ), .C1(\U8_U3_U1_n_0[0] ), 
      .C2(\U8_U3_U1_n_0[2] ), .ZN());
  XNOR2_X1_LVT U8_U3_U0_i_0_0 (.A(1'b0), .B(U8_C[3]), .ZN(
      \U8_U3_U0_DC_output[1] [15]));
  XNOR2_X1_LVT U8_U3_U0_i_0_1 (.A(\U8_U3_U0_DC_output[1] [15]), .B(1'b0), .ZN());
  INV_X1_LVT U9_U0_U0_U1_i_0_0 (.A(ci), .ZN(\U9_U0_U0_U1_n_0[0] ));
  INV_X1_LVT U9_U0_U0_U1_i_0_1 (.A(1'bz), .ZN(\U9_U0_U0_U1_n_0[1] ));
  INV_X1_LVT U9_U0_U0_U1_i_0_2 (.A(U9_C[0]), .ZN(\U9_U0_U0_U1_n_0[2] ));
  OAI222_X1_LVT U9_U0_U0_U1_i_0_3 (.A1(\U9_U0_U0_U1_n_0[0] ), .A2(
      \U9_U0_U0_U1_n_0[1] ), .B1(\U9_U0_U0_U1_n_0[1] ), .B2(\U9_U0_U0_U1_n_0[2] ), 
      .C1(\U9_U0_U0_U1_n_0[0] ), .C2(\U9_U0_U0_U1_n_0[2] ), .ZN(U9_U0_C[1]));
  XNOR2_X1_LVT U9_U0_U0_U0_i_0_0 (.A(ci), .B(U9_C[0]), .ZN(
      \U9_U0_U0_U0_DC_output[1] [15]));
  XNOR2_X1_LVT U9_U0_U0_U0_i_0_1 (.A(\U9_U0_U0_U0_DC_output[1] [15]), .B(1'bz), 
      .ZN());
  INV_X1_LVT U9_U0_U1_U1_i_0_0 (.A(ci), .ZN(\U9_U0_U1_U1_n_0[0] ));
  INV_X1_LVT U9_U0_U1_U1_i_0_1 (.A(1'b0), .ZN(\U9_U0_U1_U1_n_0[1] ));
  INV_X1_LVT U9_U0_U1_U1_i_0_2 (.A(U9_U0_C[1]), .ZN(\U9_U0_U1_U1_n_0[2] ));
  OAI222_X1_LVT U9_U0_U1_U1_i_0_3 (.A1(\U9_U0_U1_U1_n_0[0] ), .A2(
      \U9_U0_U1_U1_n_0[1] ), .B1(\U9_U0_U1_U1_n_0[1] ), .B2(\U9_U0_U1_U1_n_0[2] ), 
      .C1(\U9_U0_U1_U1_n_0[0] ), .C2(\U9_U0_U1_U1_n_0[2] ), .ZN(U9_U0_C[2]));
  XNOR2_X1_LVT U9_U0_U1_U0_i_0_0 (.A(ci), .B(U9_U0_C[1]), .ZN(
      \U9_U0_U1_U0_DC_output[1] [15]));
  XNOR2_X1_LVT U9_U0_U1_U0_i_0_1 (.A(\U9_U0_U1_U0_DC_output[1] [15]), .B(1'b0), 
      .ZN());
  INV_X1_LVT U9_U0_U2_U1_i_0_0 (.A(1'b0), .ZN(\U9_U0_U2_U1_n_0[0] ));
  INV_X1_LVT U9_U0_U2_U1_i_0_1 (.A(1'bx), .ZN(\U9_U0_U2_U1_n_0[1] ));
  INV_X1_LVT U9_U0_U2_U1_i_0_2 (.A(U9_U0_C[2]), .ZN(\U9_U0_U2_U1_n_0[2] ));
  OAI222_X1_LVT U9_U0_U2_U1_i_0_3 (.A1(\U9_U0_U2_U1_n_0[0] ), .A2(
      \U9_U0_U2_U1_n_0[1] ), .B1(\U9_U0_U2_U1_n_0[1] ), .B2(\U9_U0_U2_U1_n_0[2] ), 
      .C1(\U9_U0_U2_U1_n_0[0] ), .C2(\U9_U0_U2_U1_n_0[2] ), .ZN(U9_U0_C[3]));
  XNOR2_X1_LVT U9_U0_U2_U0_i_0_0 (.A(1'b0), .B(U9_U0_C[2]), .ZN(
      \U9_U0_U2_U0_DC_output[1] [15]));
  XNOR2_X1_LVT U9_U0_U2_U0_i_0_1 (.A(\U9_U0_U2_U0_DC_output[1] [15]), .B(1'bx), 
      .ZN());
  INV_X1_LVT U9_U0_U3_U1_i_0_0 (.A(1'b0), .ZN(\U9_U0_U3_U1_n_0[0] ));
  INV_X1_LVT U9_U0_U3_U1_i_0_1 (.A(1'b1), .ZN(\U9_U0_U3_U1_n_0[1] ));
  INV_X1_LVT U9_U0_U3_U1_i_0_2 (.A(U9_U0_C[3]), .ZN(\U9_U0_U3_U1_n_0[2] ));
  OAI222_X1_LVT U9_U0_U3_U1_i_0_3 (.A1(\U9_U0_U3_U1_n_0[0] ), .A2(
      \U9_U0_U3_U1_n_0[1] ), .B1(\U9_U0_U3_U1_n_0[1] ), .B2(\U9_U0_U3_U1_n_0[2] ), 
      .C1(\U9_U0_U3_U1_n_0[0] ), .C2(\U9_U0_U3_U1_n_0[2] ), .ZN(U9_C[1]));
  XNOR2_X1_LVT U9_U0_U3_U0_i_0_0 (.A(1'b0), .B(U9_U0_C[3]), .ZN(
      \U9_U0_U3_U0_DC_output[1] [15]));
  XNOR2_X1_LVT U9_U0_U3_U0_i_0_1 (.A(\U9_U0_U3_U0_DC_output[1] [15]), .B(1'b1), 
      .ZN());
  INV_X1_LVT U9_U1_U0_U1_i_0_0 (.A(ci), .ZN(\U9_U1_U0_U1_n_0[0] ));
  INV_X1_LVT U9_U1_U0_U1_i_0_1 (.A(1'bz), .ZN(\U9_U1_U0_U1_n_0[1] ));
  INV_X1_LVT U9_U1_U0_U1_i_0_2 (.A(U9_C[1]), .ZN(\U9_U1_U0_U1_n_0[2] ));
  OAI222_X1_LVT U9_U1_U0_U1_i_0_3 (.A1(\U9_U1_U0_U1_n_0[0] ), .A2(
      \U9_U1_U0_U1_n_0[1] ), .B1(\U9_U1_U0_U1_n_0[1] ), .B2(\U9_U1_U0_U1_n_0[2] ), 
      .C1(\U9_U1_U0_U1_n_0[0] ), .C2(\U9_U1_U0_U1_n_0[2] ), .ZN(U9_U1_C[1]));
  XNOR2_X1_LVT U9_U1_U0_U0_i_0_0 (.A(ci), .B(U9_C[1]), .ZN(
      \U9_U1_U0_U0_DC_output[1] [15]));
  XNOR2_X1_LVT U9_U1_U0_U0_i_0_1 (.A(\U9_U1_U0_U0_DC_output[1] [15]), .B(1'bz), 
      .ZN());
  INV_X1_LVT U9_U1_U1_U1_i_0_0 (.A(ci), .ZN(\U9_U1_U1_U1_n_0[0] ));
  INV_X1_LVT U9_U1_U1_U1_i_0_1 (.A(1'bx), .ZN(\U9_U1_U1_U1_n_0[1] ));
  INV_X1_LVT U9_U1_U1_U1_i_0_2 (.A(U9_U1_C[1]), .ZN(\U9_U1_U1_U1_n_0[2] ));
  OAI222_X1_LVT U9_U1_U1_U1_i_0_3 (.A1(\U9_U1_U1_U1_n_0[0] ), .A2(
      \U9_U1_U1_U1_n_0[1] ), .B1(\U9_U1_U1_U1_n_0[1] ), .B2(\U9_U1_U1_U1_n_0[2] ), 
      .C1(\U9_U1_U1_U1_n_0[0] ), .C2(\U9_U1_U1_U1_n_0[2] ), .ZN(U9_U1_C[2]));
  XNOR2_X1_LVT U9_U1_U1_U0_i_0_0 (.A(ci), .B(U9_U1_C[1]), .ZN(
      \U9_U1_U1_U0_DC_output[1] [15]));
  XNOR2_X1_LVT U9_U1_U1_U0_i_0_1 (.A(\U9_U1_U1_U0_DC_output[1] [15]), .B(1'bx), 
      .ZN());
  INV_X1_LVT U9_U1_U2_U1_i_0_0 (.A(1'b0), .ZN(\U9_U1_U2_U1_n_0[0] ));
  INV_X1_LVT U9_U1_U2_U1_i_0_1 (.A(1'b1), .ZN(\U9_U1_U2_U1_n_0[1] ));
  INV_X1_LVT U9_U1_U2_U1_i_0_2 (.A(U9_U1_C[2]), .ZN(\U9_U1_U2_U1_n_0[2] ));
  OAI222_X1_LVT U9_U1_U2_U1_i_0_3 (.A1(\U9_U1_U2_U1_n_0[0] ), .A2(
      \U9_U1_U2_U1_n_0[1] ), .B1(\U9_U1_U2_U1_n_0[1] ), .B2(\U9_U1_U2_U1_n_0[2] ), 
      .C1(\U9_U1_U2_U1_n_0[0] ), .C2(\U9_U1_U2_U1_n_0[2] ), .ZN(U9_U1_C[3]));
  XNOR2_X1_LVT U9_U1_U2_U0_i_0_0 (.A(1'b0), .B(U9_U1_C[2]), .ZN(
      \U9_U1_U2_U0_DC_output[1] [15]));
  XNOR2_X1_LVT U9_U1_U2_U0_i_0_1 (.A(\U9_U1_U2_U0_DC_output[1] [15]), .B(1'b1), 
      .ZN());
  INV_X1_LVT U9_U1_U3_U1_i_0_0 (.A(1'b0), .ZN(\U9_U1_U3_U1_n_0[0] ));
  INV_X1_LVT U9_U1_U3_U1_i_0_1 (.A(1'b0), .ZN(\U9_U1_U3_U1_n_0[1] ));
  INV_X1_LVT U9_U1_U3_U1_i_0_2 (.A(U9_U1_C[3]), .ZN(\U9_U1_U3_U1_n_0[2] ));
  OAI222_X1_LVT U9_U1_U3_U1_i_0_3 (.A1(\U9_U1_U3_U1_n_0[0] ), .A2(
      \U9_U1_U3_U1_n_0[1] ), .B1(\U9_U1_U3_U1_n_0[1] ), .B2(\U9_U1_U3_U1_n_0[2] ), 
      .C1(\U9_U1_U3_U1_n_0[0] ), .C2(\U9_U1_U3_U1_n_0[2] ), .ZN(U9_C[2]));
  XNOR2_X1_LVT U9_U1_U3_U0_i_0_0 (.A(1'b0), .B(U9_U1_C[3]), .ZN(
      \U9_U1_U3_U0_DC_output[1] [15]));
  XNOR2_X1_LVT U9_U1_U3_U0_i_0_1 (.A(\U9_U1_U3_U0_DC_output[1] [15]), .B(1'b0), 
      .ZN());
  INV_X1_LVT U9_U2_U0_U1_i_0_0 (.A(ci), .ZN(\U9_U2_U0_U1_n_0[0] ));
  INV_X1_LVT U9_U2_U0_U1_i_0_1 (.A(1'bx), .ZN(\U9_U2_U0_U1_n_0[1] ));
  INV_X1_LVT U9_U2_U0_U1_i_0_2 (.A(U9_C[2]), .ZN(\U9_U2_U0_U1_n_0[2] ));
  OAI222_X1_LVT U9_U2_U0_U1_i_0_3 (.A1(\U9_U2_U0_U1_n_0[0] ), .A2(
      \U9_U2_U0_U1_n_0[1] ), .B1(\U9_U2_U0_U1_n_0[1] ), .B2(\U9_U2_U0_U1_n_0[2] ), 
      .C1(\U9_U2_U0_U1_n_0[0] ), .C2(\U9_U2_U0_U1_n_0[2] ), .ZN(U9_U2_C[1]));
  XNOR2_X1_LVT U9_U2_U0_U0_i_0_0 (.A(ci), .B(U9_C[2]), .ZN(
      \U9_U2_U0_U0_DC_output[1] [15]));
  XNOR2_X1_LVT U9_U2_U0_U0_i_0_1 (.A(\U9_U2_U0_U0_DC_output[1] [15]), .B(1'bx), 
      .ZN());
  INV_X1_LVT U9_U2_U1_U1_i_0_0 (.A(ci), .ZN(\U9_U2_U1_U1_n_0[0] ));
  INV_X1_LVT U9_U2_U1_U1_i_0_1 (.A(ci), .ZN(\U9_U2_U1_U1_n_0[1] ));
  INV_X1_LVT U9_U2_U1_U1_i_0_2 (.A(U9_U2_C[1]), .ZN(\U9_U2_U1_U1_n_0[2] ));
  OAI222_X1_LVT U9_U2_U1_U1_i_0_3 (.A1(\U9_U2_U1_U1_n_0[0] ), .A2(
      \U9_U2_U1_U1_n_0[1] ), .B1(\U9_U2_U1_U1_n_0[1] ), .B2(\U9_U2_U1_U1_n_0[2] ), 
      .C1(\U9_U2_U1_U1_n_0[0] ), .C2(\U9_U2_U1_U1_n_0[2] ), .ZN(U9_U2_C[2]));
  XNOR2_X1_LVT U9_U2_U1_U0_i_0_0 (.A(ci), .B(U9_U2_C[1]), .ZN(
      \U9_U2_U1_U0_DC_output[1] [15]));
  XNOR2_X1_LVT U9_U2_U1_U0_i_0_1 (.A(\U9_U2_U1_U0_DC_output[1] [15]), .B(ci), 
      .ZN());
  INV_X1_LVT U9_U2_U2_U1_i_0_0 (.A(1'b0), .ZN(\U9_U2_U2_U1_n_0[0] ));
  INV_X1_LVT U9_U2_U2_U1_i_0_1 (.A(1'bz), .ZN(\U9_U2_U2_U1_n_0[1] ));
  INV_X1_LVT U9_U2_U2_U1_i_0_2 (.A(U9_U2_C[2]), .ZN(\U9_U2_U2_U1_n_0[2] ));
  OAI222_X1_LVT U9_U2_U2_U1_i_0_3 (.A1(\U9_U2_U2_U1_n_0[0] ), .A2(
      \U9_U2_U2_U1_n_0[1] ), .B1(\U9_U2_U2_U1_n_0[1] ), .B2(\U9_U2_U2_U1_n_0[2] ), 
      .C1(\U9_U2_U2_U1_n_0[0] ), .C2(\U9_U2_U2_U1_n_0[2] ), .ZN(U9_U2_C[3]));
  XNOR2_X1_LVT U9_U2_U2_U0_i_0_0 (.A(1'b0), .B(U9_U2_C[2]), .ZN(
      \U9_U2_U2_U0_DC_output[1] [15]));
  XNOR2_X1_LVT U9_U2_U2_U0_i_0_1 (.A(\U9_U2_U2_U0_DC_output[1] [15]), .B(1'bz), 
      .ZN());
  INV_X1_LVT U9_U2_U3_U1_i_0_0 (.A(1'b0), .ZN(\U9_U2_U3_U1_n_0[0] ));
  INV_X1_LVT U9_U2_U3_U1_i_0_1 (.A(1'b0), .ZN(\U9_U2_U3_U1_n_0[1] ));
  INV_X1_LVT U9_U2_U3_U1_i_0_2 (.A(U9_U2_C[3]), .ZN(\U9_U2_U3_U1_n_0[2] ));
  OAI222_X1_LVT U9_U2_U3_U1_i_0_3 (.A1(\U9_U2_U3_U1_n_0[0] ), .A2(
      \U9_U2_U3_U1_n_0[1] ), .B1(\U9_U2_U3_U1_n_0[1] ), .B2(\U9_U2_U3_U1_n_0[2] ), 
      .C1(\U9_U2_U3_U1_n_0[0] ), .C2(\U9_U2_U3_U1_n_0[2] ), .ZN(U9_c_no_defined));
  XNOR2_X1_LVT U9_U2_U3_U0_i_0_0 (.A(1'b0), .B(U9_U2_C[3]), .ZN(
      \U9_U2_U3_U0_DC_output[1] [15]));
  XNOR2_X1_LVT U9_U2_U3_U0_i_0_1 (.A(\U9_U2_U3_U0_DC_output[1] [15]), .B(1'b0), 
      .ZN());
endmodule

