module has_bigger_constant_value(B,A,C);
   inout [120:0]B;
   input [120:0]A;
   output [333:0]C;
   wire [63:0]slongv;
   wire [127:0]longv;
   wire [255:0]llongv;
  assign slongv[63] = 1'b0;
  assign slongv[62] = 1'b0;
  assign slongv[61] = 1'b0;
  assign slongv[60] = 1'b0;
  assign slongv[59] = 1'b0;
  assign slongv[58] = 1'b0;
  assign slongv[57] = 1'b0;
  assign slongv[56] = 1'b0;
  assign slongv[55] = 1'b0;
  assign slongv[54] = 1'b0;
  assign slongv[53] = 1'b0;
  assign slongv[52] = 1'b0;
  assign slongv[51] = 1'b0;
  assign slongv[50] = 1'b0;
  assign slongv[49] = 1'b0;
  assign slongv[48] = 1'b0;
  assign slongv[47] = 1'b0;
  assign slongv[46] = 1'b0;
  assign slongv[45] = 1'b0;
  assign slongv[44] = 1'b0;
  assign slongv[43] = 1'b0;
  assign slongv[42] = 1'b0;
  assign slongv[41] = 1'b0;
  assign slongv[40] = 1'b0;
  assign slongv[39] = 1'b0;
  assign slongv[38] = 1'b0;
  assign slongv[37] = 1'b0;
  assign slongv[36] = 1'b0;
  assign slongv[35] = 1'b0;
  assign slongv[34] = 1'b0;
  assign slongv[33] = 1'b1;
  assign slongv[32] = 1'b0;
  assign slongv[31] = 1'b0;
  assign slongv[30] = 1'b0;
  assign slongv[29] = 1'b0;
  assign slongv[28] = 1'b0;
  assign slongv[27] = 1'b0;
  assign slongv[26] = 1'b0;
  assign slongv[25] = 1'b0;
  assign slongv[24] = 1'b0;
  assign slongv[23] = 1'b0;
  assign slongv[22] = 1'b0;
  assign slongv[21] = 1'b0;
  assign slongv[20] = 1'b0;
  assign slongv[19] = 1'b0;
  assign slongv[18] = 1'b0;
  assign slongv[17] = 1'b0;
  assign slongv[16] = 1'b0;
  assign slongv[15] = 1'b0;
  assign slongv[14] = 1'b0;
  assign slongv[13] = 1'b0;
  assign slongv[12] = 1'b0;
  assign slongv[11] = 1'b0;
  assign slongv[10] = 1'b0;
  assign slongv[9] = 1'b0;
  assign slongv[8] = 1'b0;
  assign slongv[7] = 1'b0;
  assign slongv[6] = 1'b0;
  assign slongv[5] = 1'b0;
  assign slongv[4] = 1'b0;
  assign slongv[3] = 1'b0;
  assign slongv[2] = 1'b0;
  assign slongv[1] = 1'b0;
  assign slongv[0] = 1'b1;
  assign longv[127] = 1'b0;
  assign longv[126] = 1'b0;
  assign longv[125] = 1'b0;
  assign longv[124] = 1'b0;
  assign longv[123] = 1'b0;
  assign longv[122] = 1'b0;
  assign longv[121] = 1'b0;
  assign longv[120] = 1'b0;
  assign longv[119] = 1'b0;
  assign longv[118] = 1'b0;
  assign longv[117] = 1'b0;
  assign longv[116] = 1'b0;
  assign longv[115] = 1'b0;
  assign longv[114] = 1'b0;
  assign longv[113] = 1'b0;
  assign longv[112] = 1'b0;
  assign longv[111] = 1'b0;
  assign longv[110] = 1'b0;
  assign longv[109] = 1'b0;
  assign longv[108] = 1'b0;
  assign longv[107] = 1'b0;
  assign longv[106] = 1'b0;
  assign longv[105] = 1'b0;
  assign longv[104] = 1'b0;
  assign longv[103] = 1'b0;
  assign longv[102] = 1'b0;
  assign longv[101] = 1'b0;
  assign longv[100] = 1'b0;
  assign longv[99] = 1'b0;
  assign longv[98] = 1'b0;
  assign longv[97] = 1'b1;
  assign longv[96] = 1'b0;
  assign longv[95] = 1'b0;
  assign longv[94] = 1'b0;
  assign longv[93] = 1'b0;
  assign longv[92] = 1'b0;
  assign longv[91] = 1'b0;
  assign longv[90] = 1'b0;
  assign longv[89] = 1'b0;
  assign longv[88] = 1'b0;
  assign longv[87] = 1'b0;
  assign longv[86] = 1'b0;
  assign longv[85] = 1'b0;
  assign longv[84] = 1'b0;
  assign longv[83] = 1'b0;
  assign longv[82] = 1'b0;
  assign longv[81] = 1'b0;
  assign longv[80] = 1'b0;
  assign longv[79] = 1'b0;
  assign longv[78] = 1'b0;
  assign longv[77] = 1'b0;
  assign longv[76] = 1'b0;
  assign longv[75] = 1'b0;
  assign longv[74] = 1'b0;
  assign longv[73] = 1'b0;
  assign longv[72] = 1'b0;
  assign longv[71] = 1'b0;
  assign longv[70] = 1'b0;
  assign longv[69] = 1'b0;
  assign longv[68] = 1'b0;
  assign longv[67] = 1'b0;
  assign longv[66] = 1'b0;
  assign longv[65] = 1'b1;
  assign longv[64] = 1'b0;
  assign longv[63] = 1'b0;
  assign longv[62] = 1'b0;
  assign longv[61] = 1'b0;
  assign longv[60] = 1'b0;
  assign longv[59] = 1'b0;
  assign longv[58] = 1'b0;
  assign longv[57] = 1'b0;
  assign longv[56] = 1'b0;
  assign longv[55] = 1'b0;
  assign longv[54] = 1'b0;
  assign longv[53] = 1'b0;
  assign longv[52] = 1'b0;
  assign longv[51] = 1'b0;
  assign longv[50] = 1'b0;
  assign longv[49] = 1'b0;
  assign longv[48] = 1'b0;
  assign longv[47] = 1'b0;
  assign longv[46] = 1'b0;
  assign longv[45] = 1'b0;
  assign longv[44] = 1'b0;
  assign longv[43] = 1'b0;
  assign longv[42] = 1'b0;
  assign longv[41] = 1'b0;
  assign longv[40] = 1'b0;
  assign longv[39] = 1'b0;
  assign longv[38] = 1'b0;
  assign longv[37] = 1'b0;
  assign longv[36] = 1'b0;
  assign longv[35] = 1'b0;
  assign longv[34] = 1'b0;
  assign longv[33] = 1'b1;
  assign longv[32] = 1'b0;
  assign longv[31] = 1'b0;
  assign longv[30] = 1'b0;
  assign longv[29] = 1'b0;
  assign longv[28] = 1'b0;
  assign longv[27] = 1'b0;
  assign longv[26] = 1'b0;
  assign longv[25] = 1'b0;
  assign longv[24] = 1'b0;
  assign longv[23] = 1'b0;
  assign longv[22] = 1'b0;
  assign longv[21] = 1'b0;
  assign longv[20] = 1'b0;
  assign longv[19] = 1'b0;
  assign longv[18] = 1'b0;
  assign longv[17] = 1'b0;
  assign longv[16] = 1'b0;
  assign longv[15] = 1'b0;
  assign longv[14] = 1'b0;
  assign longv[13] = 1'b0;
  assign longv[12] = 1'b0;
  assign longv[11] = 1'b0;
  assign longv[10] = 1'b0;
  assign longv[9] = 1'b0;
  assign longv[8] = 1'b0;
  assign longv[7] = 1'b0;
  assign longv[6] = 1'b0;
  assign longv[5] = 1'b0;
  assign longv[4] = 1'b0;
  assign longv[3] = 1'b0;
  assign longv[2] = 1'b0;
  assign longv[1] = 1'b0;
  assign longv[0] = 1'b1;
  assign llongv[255] = 1'b0;
  assign llongv[254] = 1'b0;
  assign llongv[253] = 1'b0;
  assign llongv[252] = 1'b0;
  assign llongv[251] = 1'b0;
  assign llongv[250] = 1'b0;
  assign llongv[249] = 1'b0;
  assign llongv[248] = 1'b0;
  assign llongv[247] = 1'b0;
  assign llongv[246] = 1'b0;
  assign llongv[245] = 1'b0;
  assign llongv[244] = 1'b0;
  assign llongv[243] = 1'b0;
  assign llongv[242] = 1'b0;
  assign llongv[241] = 1'b0;
  assign llongv[240] = 1'b0;
  assign llongv[239] = 1'b0;
  assign llongv[238] = 1'b0;
  assign llongv[237] = 1'b0;
  assign llongv[236] = 1'b0;
  assign llongv[235] = 1'b0;
  assign llongv[234] = 1'b0;
  assign llongv[233] = 1'b0;
  assign llongv[232] = 1'b0;
  assign llongv[231] = 1'b0;
  assign llongv[230] = 1'b0;
  assign llongv[229] = 1'b0;
  assign llongv[228] = 1'b0;
  assign llongv[227] = 1'b0;
  assign llongv[226] = 1'b0;
  assign llongv[225] = 1'b1;
  assign llongv[224] = 1'b0;
  assign llongv[223] = 1'b0;
  assign llongv[222] = 1'b0;
  assign llongv[221] = 1'b0;
  assign llongv[220] = 1'b0;
  assign llongv[219] = 1'b0;
  assign llongv[218] = 1'b0;
  assign llongv[217] = 1'b0;
  assign llongv[216] = 1'b0;
  assign llongv[215] = 1'b0;
  assign llongv[214] = 1'b0;
  assign llongv[213] = 1'b0;
  assign llongv[212] = 1'b0;
  assign llongv[211] = 1'b0;
  assign llongv[210] = 1'b0;
  assign llongv[209] = 1'b0;
  assign llongv[208] = 1'b0;
  assign llongv[207] = 1'b0;
  assign llongv[206] = 1'b0;
  assign llongv[205] = 1'b0;
  assign llongv[204] = 1'b0;
  assign llongv[203] = 1'b0;
  assign llongv[202] = 1'b0;
  assign llongv[201] = 1'b0;
  assign llongv[200] = 1'b0;
  assign llongv[199] = 1'b0;
  assign llongv[198] = 1'b0;
  assign llongv[197] = 1'b0;
  assign llongv[196] = 1'b0;
  assign llongv[195] = 1'b0;
  assign llongv[194] = 1'b0;
  assign llongv[193] = 1'b0;
  assign llongv[192] = 1'b1;
  assign llongv[191] = 1'b0;
  assign llongv[190] = 1'b0;
  assign llongv[189] = 1'b0;
  assign llongv[188] = 1'b0;
  assign llongv[187] = 1'b0;
  assign llongv[186] = 1'b0;
  assign llongv[185] = 1'b0;
  assign llongv[184] = 1'b0;
  assign llongv[183] = 1'b0;
  assign llongv[182] = 1'b0;
  assign llongv[181] = 1'b0;
  assign llongv[180] = 1'b0;
  assign llongv[179] = 1'b0;
  assign llongv[178] = 1'b0;
  assign llongv[177] = 1'b0;
  assign llongv[176] = 1'b0;
  assign llongv[175] = 1'b0;
  assign llongv[174] = 1'b0;
  assign llongv[173] = 1'b0;
  assign llongv[172] = 1'b0;
  assign llongv[171] = 1'b0;
  assign llongv[170] = 1'b0;
  assign llongv[169] = 1'b0;
  assign llongv[168] = 1'b0;
  assign llongv[167] = 1'b0;
  assign llongv[166] = 1'b0;
  assign llongv[165] = 1'b0;
  assign llongv[164] = 1'b0;
  assign llongv[163] = 1'b0;
  assign llongv[162] = 1'b0;
  assign llongv[161] = 1'b1;
  assign llongv[160] = 1'b0;
  assign llongv[159] = 1'b0;
  assign llongv[158] = 1'b0;
  assign llongv[157] = 1'b0;
  assign llongv[156] = 1'b0;
  assign llongv[155] = 1'b0;
  assign llongv[154] = 1'b0;
  assign llongv[153] = 1'b0;
  assign llongv[152] = 1'b0;
  assign llongv[151] = 1'b0;
  assign llongv[150] = 1'b0;
  assign llongv[149] = 1'b0;
  assign llongv[148] = 1'b0;
  assign llongv[147] = 1'b0;
  assign llongv[146] = 1'b0;
  assign llongv[145] = 1'b0;
  assign llongv[144] = 1'b0;
  assign llongv[143] = 1'b0;
  assign llongv[142] = 1'b0;
  assign llongv[141] = 1'b0;
  assign llongv[140] = 1'b0;
  assign llongv[139] = 1'b0;
  assign llongv[138] = 1'b0;
  assign llongv[137] = 1'b0;
  assign llongv[136] = 1'b0;
  assign llongv[135] = 1'b0;
  assign llongv[134] = 1'b0;
  assign llongv[133] = 1'b0;
  assign llongv[132] = 1'b0;
  assign llongv[131] = 1'b0;
  assign llongv[130] = 1'b0;
  assign llongv[129] = 1'b1;
  assign llongv[128] = 1'b0;
  assign llongv[127] = 1'b0;
  assign llongv[126] = 1'b0;
  assign llongv[125] = 1'b0;
  assign llongv[124] = 1'b0;
  assign llongv[123] = 1'b0;
  assign llongv[122] = 1'b0;
  assign llongv[121] = 1'b0;
  assign llongv[120] = 1'b0;
  assign llongv[119] = 1'b0;
  assign llongv[118] = 1'b0;
  assign llongv[117] = 1'b0;
  assign llongv[116] = 1'b0;
  assign llongv[115] = 1'b0;
  assign llongv[114] = 1'b0;
  assign llongv[113] = 1'b0;
  assign llongv[112] = 1'b0;
  assign llongv[111] = 1'b0;
  assign llongv[110] = 1'b0;
  assign llongv[109] = 1'b0;
  assign llongv[108] = 1'b0;
  assign llongv[107] = 1'b0;
  assign llongv[106] = 1'b0;
  assign llongv[105] = 1'b0;
  assign llongv[104] = 1'b0;
  assign llongv[103] = 1'b0;
  assign llongv[102] = 1'b0;
  assign llongv[101] = 1'b0;
  assign llongv[100] = 1'b0;
  assign llongv[99] = 1'b0;
  assign llongv[98] = 1'b0;
  assign llongv[97] = 1'b1;
  assign llongv[96] = 1'b0;
  assign llongv[95] = 1'b0;
  assign llongv[94] = 1'b0;
  assign llongv[93] = 1'b0;
  assign llongv[92] = 1'b0;
  assign llongv[91] = 1'b0;
  assign llongv[90] = 1'b0;
  assign llongv[89] = 1'b0;
  assign llongv[88] = 1'b0;
  assign llongv[87] = 1'b0;
  assign llongv[86] = 1'b0;
  assign llongv[85] = 1'b0;
  assign llongv[84] = 1'b0;
  assign llongv[83] = 1'b0;
  assign llongv[82] = 1'b0;
  assign llongv[81] = 1'b0;
  assign llongv[80] = 1'b0;
  assign llongv[79] = 1'b0;
  assign llongv[78] = 1'b0;
  assign llongv[77] = 1'b0;
  assign llongv[76] = 1'b0;
  assign llongv[75] = 1'b0;
  assign llongv[74] = 1'b0;
  assign llongv[73] = 1'b0;
  assign llongv[72] = 1'b0;
  assign llongv[71] = 1'b0;
  assign llongv[70] = 1'b0;
  assign llongv[69] = 1'b0;
  assign llongv[68] = 1'b0;
  assign llongv[67] = 1'b0;
  assign llongv[66] = 1'b0;
  assign llongv[65] = 1'b0;
  assign llongv[64] = 1'b1;
  assign llongv[63] = 1'b0;
  assign llongv[62] = 1'b0;
  assign llongv[61] = 1'b0;
  assign llongv[60] = 1'b0;
  assign llongv[59] = 1'b0;
  assign llongv[58] = 1'b0;
  assign llongv[57] = 1'b0;
  assign llongv[56] = 1'b0;
  assign llongv[55] = 1'b0;
  assign llongv[54] = 1'b0;
  assign llongv[53] = 1'b0;
  assign llongv[52] = 1'b0;
  assign llongv[51] = 1'b0;
  assign llongv[50] = 1'b0;
  assign llongv[49] = 1'b0;
  assign llongv[48] = 1'b0;
  assign llongv[47] = 1'b0;
  assign llongv[46] = 1'b0;
  assign llongv[45] = 1'b0;
  assign llongv[44] = 1'b0;
  assign llongv[43] = 1'b0;
  assign llongv[42] = 1'b0;
  assign llongv[41] = 1'b0;
  assign llongv[40] = 1'b0;
  assign llongv[39] = 1'b0;
  assign llongv[38] = 1'b0;
  assign llongv[37] = 1'b0;
  assign llongv[36] = 1'b0;
  assign llongv[35] = 1'b0;
  assign llongv[34] = 1'b0;
  assign llongv[33] = 1'b1;
  assign llongv[32] = 1'b0;
  assign llongv[31] = 1'b0;
  assign llongv[30] = 1'b0;
  assign llongv[29] = 1'b0;
  assign llongv[28] = 1'b0;
  assign llongv[27] = 1'b0;
  assign llongv[26] = 1'b0;
  assign llongv[25] = 1'b0;
  assign llongv[24] = 1'b0;
  assign llongv[23] = 1'b0;
  assign llongv[22] = 1'b0;
  assign llongv[21] = 1'b0;
  assign llongv[20] = 1'b0;
  assign llongv[19] = 1'b0;
  assign llongv[18] = 1'b0;
  assign llongv[17] = 1'b0;
  assign llongv[16] = 1'b0;
  assign llongv[15] = 1'b0;
  assign llongv[14] = 1'b0;
  assign llongv[13] = 1'b0;
  assign llongv[12] = 1'b0;
  assign llongv[11] = 1'b0;
  assign llongv[10] = 1'b0;
  assign llongv[9] = 1'b0;
  assign llongv[8] = 1'b0;
  assign llongv[7] = 1'b0;
  assign llongv[6] = 1'b0;
  assign llongv[5] = 1'b0;
  assign llongv[4] = 1'b0;
  assign llongv[3] = 1'b0;
  assign llongv[2] = 1'b0;
  assign llongv[1] = 1'b0;
  assign llongv[0] = 1'b1;
  assign C[64] = B[64];
  assign C[63] = B[63];
  assign C[62] = B[62];
  assign C[61] = B[61];
  assign C[60] = B[60];
  assign C[59] = B[59];
  assign C[58] = B[58];
  assign C[57] = B[57];
  assign C[56] = B[56];
  assign C[55] = B[55];
  assign C[54] = B[54];
  assign C[53] = B[53];
  assign C[52] = B[52];
  assign C[51] = B[51];
  assign C[50] = B[50];
  assign C[49] = B[49];
  assign C[48] = B[48];
  assign C[47] = B[47];
  assign C[46] = B[46];
  assign C[45] = B[45];
  assign C[44] = B[44];
  assign C[43] = B[43];
  assign C[42] = B[42];
  assign C[41] = B[41];
  assign C[40] = B[40];
  assign C[39] = B[39];
  assign C[38] = B[38];
  assign C[37] = B[37];
  assign C[36] = B[36];
  assign C[105] = B[105];
  assign C[104] = B[104];
  assign C[103] = B[103];
  assign C[102] = B[102];
  assign C[101] = B[101];
  assign C[100] = B[100];
  assign C[99] = B[99];
  assign C[98] = B[98];
  assign C[97] = B[97];
  assign C[96] = B[96];
  assign C[95] = B[95];
  assign C[94] = B[94];
  assign C[93] = B[93];
  assign C[92] = B[92];
  assign C[91] = B[91];
  assign C[90] = B[90];
  assign C[89] = B[89];
  assign C[88] = B[88];
  assign C[87] = B[87];
  assign C[86] = B[86];
  assign C[85] = B[85];
  assign C[84] = B[84];
  assign C[83] = B[83];
  assign C[82] = B[82];
  assign C[81] = B[81];
  assign C[80] = B[80];
  assign C[79] = B[79];
  assign C[78] = B[78];
  assign C[77] = B[77];
  assign C[170] = longv[105];
  assign C[169] = longv[104];
  assign C[168] = longv[103];
  assign C[167] = longv[102];
  assign C[166] = longv[101];
  assign C[165] = longv[100];
  assign C[164] = longv[99];
  assign C[163] = longv[98];
  assign C[162] = longv[97];
  assign C[161] = longv[96];
  assign C[160] = longv[95];
  assign C[159] = longv[94];
  assign C[158] = longv[93];
  assign C[157] = longv[92];
  assign C[156] = longv[91];
  assign C[155] = longv[90];
  assign C[154] = longv[89];
  assign C[153] = longv[88];
  assign C[152] = longv[87];
  assign C[151] = longv[86];
  assign C[150] = longv[85];
  assign C[149] = longv[84];
  assign C[148] = longv[83];
  assign C[147] = longv[82];
  assign C[146] = longv[81];
  assign C[145] = longv[80];
  assign C[144] = longv[79];
  assign C[143] = longv[78];
  assign C[142] = longv[77];
  INV_X1_LVT U1/U1/i_0_0 (.A(A[0]), .ZN(C[0]));
  INV_X1_LVT U1/U1/i_0_1 (.A(B[0]), .ZN(C[1]));
  INV_X1_LVT U1/U1/i_0_2 (.A(B[1]), .ZN(C[2]));
  OAI222_X1_LVT U1/U1/i_0_3 (.A1(A[1]), .A2(A[2]), .B1(B[1]), .B2(B[2]), .C1(
      A[3]), .C2(B[3]), .ZN(C[3]));
  INV_X1_LVT U1/U1/i_1_0 (.A(A[4]), .ZN(C[4]));
  INV_X1_LVT U1/U1/i_1_1 (.A(B[4]), .ZN(C[5]));
  INV_X1_LVT U1/U1/i_1_2 (.A(B[5]), .ZN(C[6]));
  OAI222_X1_LVT U1/U1/i_1_3 (.A1(A[5]), .A2(A[6]), .B1(B[5]), .B2(B[6]), .C1(
      A[7]), .C2(B[7]), .ZN(C[7]));
  INV_X1_LVT U1/U1/i_2_0 (.A(A[8]), .ZN(C[8]));
  INV_X1_LVT U1/U1/i_2_1 (.A(B[8]), .ZN(C[9]));
  INV_X1_LVT U1/U1/i_2_2 (.A(B[9]), .ZN(C[10]));
  OAI222_X1_LVT U1/U1/i_2_3 (.A1(A[9]), .A2(A[10]), .B1(B[9]), .B2(B[10]), .C1(
      A[11]), .C2(B[11]), .ZN(C[11]));
  INV_X1_LVT U1/U2/i_0_0 (.A(A[12]), .ZN(C[12]));
  INV_X1_LVT U1/U2/i_0_1 (.A(B[12]), .ZN(C[13]));
  INV_X1_LVT U1/U2/i_0_2 (.A(B[13]), .ZN(C[14]));
  OAI222_X1_LVT U1/U2/i_0_3 (.A1(A[13]), .A2(A[14]), .B1(B[13]), .B2(B[14]), .C1(
      A[15]), .C2(B[15]), .ZN(C[15]));
  INV_X1_LVT U1/U2/i_1_0 (.A(A[16]), .ZN(C[16]));
  INV_X1_LVT U1/U2/i_1_1 (.A(B[16]), .ZN(C[17]));
  INV_X1_LVT U1/U2/i_1_2 (.A(B[17]), .ZN(C[18]));
  OAI222_X1_LVT U1/U2/i_1_3 (.A1(A[17]), .A2(A[18]), .B1(B[17]), .B2(B[18]), .C1(
      A[19]), .C2(B[19]), .ZN(C[19]));
  INV_X1_LVT U1/U2/i_2_0 (.A(A[20]), .ZN(C[20]));
  INV_X1_LVT U1/U2/i_2_1 (.A(B[20]), .ZN(C[21]));
  INV_X1_LVT U1/U2/i_2_2 (.A(B[21]), .ZN(C[22]));
  OAI222_X1_LVT U1/U2/i_2_3 (.A1(A[21]), .A2(A[22]), .B1(B[21]), .B2(B[22]), .C1(
      A[23]), .C2(B[23]), .ZN(C[23]));
  INV_X1_LVT U1/U3/i_0_0 (.A(A[24]), .ZN(C[24]));
  INV_X1_LVT U1/U3/i_0_1 (.A(B[24]), .ZN(C[25]));
  INV_X1_LVT U1/U3/i_0_2 (.A(B[25]), .ZN(C[26]));
  OAI222_X1_LVT U1/U3/i_0_3 (.A1(A[25]), .A2(A[26]), .B1(B[25]), .B2(B[26]), .C1(
      A[27]), .C2(B[27]), .ZN(C[27]));
  INV_X1_LVT U1/U3/i_1_0 (.A(A[28]), .ZN(C[28]));
  INV_X1_LVT U1/U3/i_1_1 (.A(B[28]), .ZN(C[29]));
  INV_X1_LVT U1/U3/i_1_2 (.A(B[29]), .ZN(C[30]));
  OAI222_X1_LVT U1/U3/i_1_3 (.A1(A[29]), .A2(A[30]), .B1(B[29]), .B2(B[30]), .C1(
      A[31]), .C2(B[31]), .ZN(C[31]));
  INV_X1_LVT U1/U3/i_2_0 (.A(A[32]), .ZN(C[32]));
  INV_X1_LVT U1/U3/i_2_1 (.A(B[32]), .ZN(C[33]));
  INV_X1_LVT U1/U3/i_2_2 (.A(B[33]), .ZN(C[34]));
  OAI222_X1_LVT U1/U3/i_2_3 (.A1(A[33]), .A2(A[34]), .B1(B[33]), .B2(B[34]), .C1(
      A[35]), .C2(B[35]), .ZN(C[35]));
  INV_X1_LVT U2/U1/i_0_0 (.A(A[41]), .ZN(C[41]));
  INV_X1_LVT U2/U1/i_0_1 (.A(B[41]), .ZN(C[42]));
  INV_X1_LVT U2/U1/i_0_2 (.A(B[42]), .ZN(C[43]));
  OAI222_X1_LVT U2/U1/i_0_3 (.A1(A[42]), .A2(A[43]), .B1(B[42]), .B2(B[43]), .C1(
      A[44]), .C2(B[44]), .ZN(C[44]));
  INV_X1_LVT U2/U1/i_1_0 (.A(A[45]), .ZN(C[45]));
  INV_X1_LVT U2/U1/i_1_1 (.A(B[45]), .ZN(C[46]));
  INV_X1_LVT U2/U1/i_1_2 (.A(B[46]), .ZN(C[47]));
  OAI222_X1_LVT U2/U1/i_1_3 (.A1(A[46]), .A2(A[47]), .B1(B[46]), .B2(B[47]), .C1(
      A[48]), .C2(B[48]), .ZN(C[48]));
  INV_X1_LVT U2/U1/i_2_0 (.A(A[49]), .ZN(C[49]));
  INV_X1_LVT U2/U1/i_2_1 (.A(B[49]), .ZN(C[50]));
  INV_X1_LVT U2/U1/i_2_2 (.A(B[50]), .ZN(C[51]));
  OAI222_X1_LVT U2/U1/i_2_3 (.A1(A[50]), .A2(A[51]), .B1(B[50]), .B2(B[51]), .C1(
      A[52]), .C2(B[52]), .ZN(C[52]));
  INV_X1_LVT U2/U2/i_0_0 (.A(A[53]), .ZN(C[53]));
  INV_X1_LVT U2/U2/i_0_1 (.A(B[53]), .ZN(C[54]));
  INV_X1_LVT U2/U2/i_0_2 (.A(B[54]), .ZN(C[55]));
  OAI222_X1_LVT U2/U2/i_0_3 (.A1(A[54]), .A2(A[55]), .B1(B[54]), .B2(B[55]), .C1(
      A[56]), .C2(B[56]), .ZN(C[56]));
  INV_X1_LVT U2/U2/i_1_0 (.A(A[57]), .ZN(C[57]));
  INV_X1_LVT U2/U2/i_1_1 (.A(B[57]), .ZN(C[58]));
  INV_X1_LVT U2/U2/i_1_2 (.A(B[58]), .ZN(C[59]));
  OAI222_X1_LVT U2/U2/i_1_3 (.A1(A[58]), .A2(A[59]), .B1(B[58]), .B2(B[59]), .C1(
      A[60]), .C2(B[60]), .ZN(C[60]));
  INV_X1_LVT U2/U2/i_2_0 (.A(A[61]), .ZN(C[61]));
  INV_X1_LVT U2/U2/i_2_1 (.A(B[61]), .ZN(C[62]));
  INV_X1_LVT U2/U2/i_2_2 (.A(B[62]), .ZN(C[63]));
  OAI222_X1_LVT U2/U2/i_2_3 (.A1(A[62]), .A2(A[63]), .B1(B[62]), .B2(B[63]), .C1(
      A[64]), .C2(B[64]), .ZN(C[64]));
  INV_X1_LVT U2/U3/i_0_0 (.A(A[65]), .ZN(C[65]));
  INV_X1_LVT U2/U3/i_0_1 (.A(B[65]), .ZN(C[66]));
  INV_X1_LVT U2/U3/i_0_2 (.A(B[66]), .ZN(C[67]));
  OAI222_X1_LVT U2/U3/i_0_3 (.A1(A[66]), .A2(A[67]), .B1(B[66]), .B2(B[67]), .C1(
      A[68]), .C2(B[68]), .ZN(C[68]));
  INV_X1_LVT U2/U3/i_1_0 (.A(A[69]), .ZN(C[69]));
  INV_X1_LVT U2/U3/i_1_1 (.A(B[69]), .ZN(C[70]));
  INV_X1_LVT U2/U3/i_1_2 (.A(B[70]), .ZN(C[71]));
  OAI222_X1_LVT U2/U3/i_1_3 (.A1(A[70]), .A2(A[71]), .B1(B[70]), .B2(B[71]), .C1(
      A[72]), .C2(B[72]), .ZN(C[72]));
  INV_X1_LVT U2/U3/i_2_0 (.A(A[73]), .ZN(C[73]));
  INV_X1_LVT U2/U3/i_2_1 (.A(B[73]), .ZN(C[74]));
  INV_X1_LVT U2/U3/i_2_2 (.A(B[74]), .ZN(C[75]));
  OAI222_X1_LVT U2/U3/i_2_3 (.A1(A[74]), .A2(A[75]), .B1(B[74]), .B2(B[75]), .C1(
      A[76]), .C2(B[76]), .ZN(C[76]));
  INV_X1_LVT U3/U1/i_0_0 (.A(1'b0), .ZN(C[106]));
  INV_X1_LVT U3/U1/i_0_1 (.A(longv[41]), .ZN(C[107]));
  INV_X1_LVT U3/U1/i_0_2 (.A(longv[42]), .ZN(C[108]));
  OAI222_X1_LVT U3/U1/i_0_3 (.A1(1'b1), .A2(1'b0), .B1(longv[42]), .B2(longv[43]), 
      .C1(1'b0), .C2(longv[44]), .ZN(C[109]));
  INV_X1_LVT U3/U1/i_1_0 (.A(1'b0), .ZN(C[110]));
  INV_X1_LVT U3/U1/i_1_1 (.A(longv[45]), .ZN(C[111]));
  INV_X1_LVT U3/U1/i_1_2 (.A(longv[46]), .ZN(C[112]));
  OAI222_X1_LVT U3/U1/i_1_3 (.A1(1'b0), .A2(1'b0), .B1(longv[46]), .B2(longv[47]), 
      .C1(1'b0), .C2(longv[48]), .ZN(C[113]));
  INV_X1_LVT U3/U1/i_2_0 (.A(1'b0), .ZN(C[114]));
  INV_X1_LVT U3/U1/i_2_1 (.A(longv[49]), .ZN(C[115]));
  INV_X1_LVT U3/U1/i_2_2 (.A(longv[50]), .ZN(C[116]));
  OAI222_X1_LVT U3/U1/i_2_3 (.A1(1'b0), .A2(1'b0), .B1(longv[50]), .B2(longv[51]), 
      .C1(1'b0), .C2(longv[52]), .ZN(C[117]));
  INV_X1_LVT U3/U2/i_0_0 (.A(1'b0), .ZN(C[118]));
  INV_X1_LVT U3/U2/i_0_1 (.A(longv[53]), .ZN(C[119]));
  INV_X1_LVT U3/U2/i_0_2 (.A(longv[54]), .ZN(C[120]));
  OAI222_X1_LVT U3/U2/i_0_3 (.A1(1'b0), .A2(1'b0), .B1(longv[54]), .B2(longv[55]), 
      .C1(1'b0), .C2(longv[56]), .ZN(C[121]));
  INV_X1_LVT U3/U2/i_1_0 (.A(1'b0), .ZN(C[122]));
  INV_X1_LVT U3/U2/i_1_1 (.A(longv[57]), .ZN(C[123]));
  INV_X1_LVT U3/U2/i_1_2 (.A(longv[58]), .ZN(C[124]));
  OAI222_X1_LVT U3/U2/i_1_3 (.A1(1'b0), .A2(1'b0), .B1(longv[58]), .B2(longv[59]), 
      .C1(1'b0), .C2(longv[60]), .ZN(C[125]));
  INV_X1_LVT U3/U2/i_2_0 (.A(1'b0), .ZN(C[126]));
  INV_X1_LVT U3/U2/i_2_1 (.A(longv[61]), .ZN(C[127]));
  INV_X1_LVT U3/U2/i_2_2 (.A(longv[62]), .ZN(C[128]));
  OAI222_X1_LVT U3/U2/i_2_3 (.A1(1'b0), .A2(1'b0), .B1(longv[62]), .B2(longv[63]), 
      .C1(1'b0), .C2(longv[64]), .ZN(C[129]));
  INV_X1_LVT U3/U3/i_0_0 (.A(1'b0), .ZN(C[130]));
  INV_X1_LVT U3/U3/i_0_1 (.A(longv[65]), .ZN(C[131]));
  INV_X1_LVT U3/U3/i_0_2 (.A(longv[66]), .ZN(C[132]));
  OAI222_X1_LVT U3/U3/i_0_3 (.A1(1'b0), .A2(1'b0), .B1(longv[66]), .B2(longv[67]), 
      .C1(1'b0), .C2(longv[68]), .ZN(C[133]));
  INV_X1_LVT U3/U3/i_1_0 (.A(1'b0), .ZN(C[134]));
  INV_X1_LVT U3/U3/i_1_1 (.A(longv[69]), .ZN(C[135]));
  INV_X1_LVT U3/U3/i_1_2 (.A(longv[70]), .ZN(C[136]));
  OAI222_X1_LVT U3/U3/i_1_3 (.A1(1'b0), .A2(1'b0), .B1(longv[70]), .B2(longv[71]), 
      .C1(1'b0), .C2(longv[72]), .ZN(C[137]));
  INV_X1_LVT U3/U3/i_2_0 (.A(1'b0), .ZN(C[138]));
  INV_X1_LVT U3/U3/i_2_1 (.A(longv[73]), .ZN(C[139]));
  INV_X1_LVT U3/U3/i_2_2 (.A(longv[74]), .ZN(C[140]));
  OAI222_X1_LVT U3/U3/i_2_3 (.A1(1'b1), .A2(1'b0), .B1(longv[74]), .B2(longv[75]), 
      .C1(1'b0), .C2(longv[76]), .ZN(C[141]));
endmodule

