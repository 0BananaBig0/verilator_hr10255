module AOTOP(a,b,c,d,e);
   input a;
   input b;
   input c;
   output d;
   output e;
  assign d = a;
endmodule

