module has_bigger_constant_value(A,B,C);
   input [120:0]A;
   inout [120:0]B;
   output [122:0]C;
   wire [63:0]slongv;
   wire [127:0]longv;
   wire [255:0]llongv;
  assign slongv[63] = 1'b0;
  assign slongv[62] = 1'b0;
  assign slongv[61] = 1'b0;
  assign slongv[60] = 1'b0;
  assign slongv[59] = 1'b0;
  assign slongv[58] = 1'b0;
  assign slongv[57] = 1'b0;
  assign slongv[56] = 1'b0;
  assign slongv[55] = 1'b0;
  assign slongv[54] = 1'b0;
  assign slongv[53] = 1'b0;
  assign slongv[52] = 1'b0;
  assign slongv[51] = 1'b0;
  assign slongv[50] = 1'b0;
  assign slongv[49] = 1'b0;
  assign slongv[48] = 1'b0;
  assign slongv[47] = 1'b0;
  assign slongv[46] = 1'b0;
  assign slongv[45] = 1'b0;
  assign slongv[44] = 1'b0;
  assign slongv[43] = 1'b0;
  assign slongv[42] = 1'b0;
  assign slongv[41] = 1'b0;
  assign slongv[40] = 1'b0;
  assign slongv[39] = 1'b0;
  assign slongv[38] = 1'b0;
  assign slongv[37] = 1'b0;
  assign slongv[36] = 1'b0;
  assign slongv[35] = 1'b0;
  assign slongv[34] = 1'b0;
  assign slongv[33] = 1'b1;
  assign slongv[32] = 1'b0;
  assign slongv[31] = 1'b0;
  assign slongv[30] = 1'b0;
  assign slongv[29] = 1'b0;
  assign slongv[28] = 1'b0;
  assign slongv[27] = 1'b0;
  assign slongv[26] = 1'b0;
  assign slongv[25] = 1'b0;
  assign slongv[24] = 1'b0;
  assign slongv[23] = 1'b0;
  assign slongv[22] = 1'b0;
  assign slongv[21] = 1'b0;
  assign slongv[20] = 1'b0;
  assign slongv[19] = 1'b0;
  assign slongv[18] = 1'b0;
  assign slongv[17] = 1'b0;
  assign slongv[16] = 1'b0;
  assign slongv[15] = 1'b0;
  assign slongv[14] = 1'b0;
  assign slongv[13] = 1'b0;
  assign slongv[12] = 1'b0;
  assign slongv[11] = 1'b0;
  assign slongv[10] = 1'b0;
  assign slongv[9] = 1'b0;
  assign slongv[8] = 1'b0;
  assign slongv[7] = 1'b0;
  assign slongv[6] = 1'b0;
  assign slongv[5] = 1'b0;
  assign slongv[4] = 1'b0;
  assign slongv[3] = 1'b0;
  assign slongv[2] = 1'b0;
  assign slongv[1] = 1'b0;
  assign slongv[0] = 1'b1;
  assign longv[127] = 1'b0;
  assign longv[126] = 1'b0;
  assign longv[125] = 1'b0;
  assign longv[124] = 1'b0;
  assign longv[123] = 1'b0;
  assign longv[122] = 1'b0;
  assign longv[121] = 1'b0;
  assign longv[120] = 1'b0;
  assign longv[119] = 1'b0;
  assign longv[118] = 1'b0;
  assign longv[117] = 1'b0;
  assign longv[116] = 1'b0;
  assign longv[115] = 1'b0;
  assign longv[114] = 1'b0;
  assign longv[113] = 1'b0;
  assign longv[112] = 1'b0;
  assign longv[111] = 1'b0;
  assign longv[110] = 1'b0;
  assign longv[109] = 1'b0;
  assign longv[108] = 1'b0;
  assign longv[107] = 1'b0;
  assign longv[106] = 1'b0;
  assign longv[105] = 1'b0;
  assign longv[104] = 1'b0;
  assign longv[103] = 1'b0;
  assign longv[102] = 1'b0;
  assign longv[101] = 1'b0;
  assign longv[100] = 1'b0;
  assign longv[99] = 1'b0;
  assign longv[98] = 1'b0;
  assign longv[97] = 1'b1;
  assign longv[96] = 1'b0;
  assign longv[95] = 1'b0;
  assign longv[94] = 1'b0;
  assign longv[93] = 1'b0;
  assign longv[92] = 1'b0;
  assign longv[91] = 1'b0;
  assign longv[90] = 1'b0;
  assign longv[89] = 1'b0;
  assign longv[88] = 1'b0;
  assign longv[87] = 1'b0;
  assign longv[86] = 1'b0;
  assign longv[85] = 1'b0;
  assign longv[84] = 1'b0;
  assign longv[83] = 1'b0;
  assign longv[82] = 1'b0;
  assign longv[81] = 1'b0;
  assign longv[80] = 1'b0;
  assign longv[79] = 1'b0;
  assign longv[78] = 1'b0;
  assign longv[77] = 1'b0;
  assign longv[76] = 1'b0;
  assign longv[75] = 1'b0;
  assign longv[74] = 1'b0;
  assign longv[73] = 1'b0;
  assign longv[72] = 1'b0;
  assign longv[71] = 1'b0;
  assign longv[70] = 1'b0;
  assign longv[69] = 1'b0;
  assign longv[68] = 1'b0;
  assign longv[67] = 1'b0;
  assign longv[66] = 1'b0;
  assign longv[65] = 1'b1;
  assign longv[64] = 1'b0;
  assign longv[63] = 1'b0;
  assign longv[62] = 1'b0;
  assign longv[61] = 1'b0;
  assign longv[60] = 1'b0;
  assign longv[59] = 1'b0;
  assign longv[58] = 1'b0;
  assign longv[57] = 1'b0;
  assign longv[56] = 1'b0;
  assign longv[55] = 1'b0;
  assign longv[54] = 1'b0;
  assign longv[53] = 1'b0;
  assign longv[52] = 1'b0;
  assign longv[51] = 1'b0;
  assign longv[50] = 1'b0;
  assign longv[49] = 1'b0;
  assign longv[48] = 1'b0;
  assign longv[47] = 1'b0;
  assign longv[46] = 1'b0;
  assign longv[45] = 1'b0;
  assign longv[44] = 1'b0;
  assign longv[43] = 1'b0;
  assign longv[42] = 1'b0;
  assign longv[41] = 1'b0;
  assign longv[40] = 1'b0;
  assign longv[39] = 1'b0;
  assign longv[38] = 1'b0;
  assign longv[37] = 1'b0;
  assign longv[36] = 1'b0;
  assign longv[35] = 1'b0;
  assign longv[34] = 1'b0;
  assign longv[33] = 1'b1;
  assign longv[32] = 1'b0;
  assign longv[31] = 1'b0;
  assign longv[30] = 1'b0;
  assign longv[29] = 1'b0;
  assign longv[28] = 1'b0;
  assign longv[27] = 1'b0;
  assign longv[26] = 1'b0;
  assign longv[25] = 1'b0;
  assign longv[24] = 1'b0;
  assign longv[23] = 1'b0;
  assign longv[22] = 1'b0;
  assign longv[21] = 1'b0;
  assign longv[20] = 1'b0;
  assign longv[19] = 1'b0;
  assign longv[18] = 1'b0;
  assign longv[17] = 1'b0;
  assign longv[16] = 1'b0;
  assign longv[15] = 1'b0;
  assign longv[14] = 1'b0;
  assign longv[13] = 1'b0;
  assign longv[12] = 1'b0;
  assign longv[11] = 1'b0;
  assign longv[10] = 1'b0;
  assign longv[9] = 1'b0;
  assign longv[8] = 1'b0;
  assign longv[7] = 1'b0;
  assign longv[6] = 1'b0;
  assign longv[5] = 1'b0;
  assign longv[4] = 1'b0;
  assign longv[3] = 1'b0;
  assign longv[2] = 1'b0;
  assign longv[1] = 1'b0;
  assign longv[0] = 1'b1;
  assign llongv[255] = 1'b0;
  assign llongv[254] = 1'b0;
  assign llongv[253] = 1'b0;
  assign llongv[252] = 1'b0;
  assign llongv[251] = 1'b0;
  assign llongv[250] = 1'b0;
  assign llongv[249] = 1'b0;
  assign llongv[248] = 1'b0;
  assign llongv[247] = 1'b0;
  assign llongv[246] = 1'b0;
  assign llongv[245] = 1'b0;
  assign llongv[244] = 1'b0;
  assign llongv[243] = 1'b0;
  assign llongv[242] = 1'b0;
  assign llongv[241] = 1'b0;
  assign llongv[240] = 1'b0;
  assign llongv[239] = 1'b0;
  assign llongv[238] = 1'b0;
  assign llongv[237] = 1'b0;
  assign llongv[236] = 1'b0;
  assign llongv[235] = 1'b0;
  assign llongv[234] = 1'b0;
  assign llongv[233] = 1'b0;
  assign llongv[232] = 1'b0;
  assign llongv[231] = 1'b0;
  assign llongv[230] = 1'b0;
  assign llongv[229] = 1'b0;
  assign llongv[228] = 1'b0;
  assign llongv[227] = 1'b0;
  assign llongv[226] = 1'b0;
  assign llongv[225] = 1'b1;
  assign llongv[224] = 1'b0;
  assign llongv[223] = 1'b0;
  assign llongv[222] = 1'b0;
  assign llongv[221] = 1'b0;
  assign llongv[220] = 1'b0;
  assign llongv[219] = 1'b0;
  assign llongv[218] = 1'b0;
  assign llongv[217] = 1'b0;
  assign llongv[216] = 1'b0;
  assign llongv[215] = 1'b0;
  assign llongv[214] = 1'b0;
  assign llongv[213] = 1'b0;
  assign llongv[212] = 1'b0;
  assign llongv[211] = 1'b0;
  assign llongv[210] = 1'b0;
  assign llongv[209] = 1'b0;
  assign llongv[208] = 1'b0;
  assign llongv[207] = 1'b0;
  assign llongv[206] = 1'b0;
  assign llongv[205] = 1'b0;
  assign llongv[204] = 1'b0;
  assign llongv[203] = 1'b0;
  assign llongv[202] = 1'b0;
  assign llongv[201] = 1'b0;
  assign llongv[200] = 1'b0;
  assign llongv[199] = 1'b0;
  assign llongv[198] = 1'b0;
  assign llongv[197] = 1'b0;
  assign llongv[196] = 1'b0;
  assign llongv[195] = 1'b0;
  assign llongv[194] = 1'b0;
  assign llongv[193] = 1'b0;
  assign llongv[192] = 1'b1;
  assign llongv[191] = 1'b0;
  assign llongv[190] = 1'b0;
  assign llongv[189] = 1'b0;
  assign llongv[188] = 1'b0;
  assign llongv[187] = 1'b0;
  assign llongv[186] = 1'b0;
  assign llongv[185] = 1'b0;
  assign llongv[184] = 1'b0;
  assign llongv[183] = 1'b0;
  assign llongv[182] = 1'b0;
  assign llongv[181] = 1'b0;
  assign llongv[180] = 1'b0;
  assign llongv[179] = 1'b0;
  assign llongv[178] = 1'b0;
  assign llongv[177] = 1'b0;
  assign llongv[176] = 1'b0;
  assign llongv[175] = 1'b0;
  assign llongv[174] = 1'b0;
  assign llongv[173] = 1'b0;
  assign llongv[172] = 1'b0;
  assign llongv[171] = 1'b0;
  assign llongv[170] = 1'b0;
  assign llongv[169] = 1'b0;
  assign llongv[168] = 1'b0;
  assign llongv[167] = 1'b0;
  assign llongv[166] = 1'b0;
  assign llongv[165] = 1'b0;
  assign llongv[164] = 1'b0;
  assign llongv[163] = 1'b0;
  assign llongv[162] = 1'b0;
  assign llongv[161] = 1'b1;
  assign llongv[160] = 1'b0;
  assign llongv[159] = 1'b0;
  assign llongv[158] = 1'b0;
  assign llongv[157] = 1'b0;
  assign llongv[156] = 1'b0;
  assign llongv[155] = 1'b0;
  assign llongv[154] = 1'b0;
  assign llongv[153] = 1'b0;
  assign llongv[152] = 1'b0;
  assign llongv[151] = 1'b0;
  assign llongv[150] = 1'b0;
  assign llongv[149] = 1'b0;
  assign llongv[148] = 1'b0;
  assign llongv[147] = 1'b0;
  assign llongv[146] = 1'b0;
  assign llongv[145] = 1'b0;
  assign llongv[144] = 1'b0;
  assign llongv[143] = 1'b0;
  assign llongv[142] = 1'b0;
  assign llongv[141] = 1'b0;
  assign llongv[140] = 1'b0;
  assign llongv[139] = 1'b0;
  assign llongv[138] = 1'b0;
  assign llongv[137] = 1'b0;
  assign llongv[136] = 1'b0;
  assign llongv[135] = 1'b0;
  assign llongv[134] = 1'b0;
  assign llongv[133] = 1'b0;
  assign llongv[132] = 1'b0;
  assign llongv[131] = 1'b0;
  assign llongv[130] = 1'b0;
  assign llongv[129] = 1'b1;
  assign llongv[128] = 1'b0;
  assign llongv[127] = 1'b0;
  assign llongv[126] = 1'b0;
  assign llongv[125] = 1'b0;
  assign llongv[124] = 1'b0;
  assign llongv[123] = 1'b0;
  assign llongv[122] = 1'b0;
  assign llongv[121] = 1'b0;
  assign llongv[120] = 1'b0;
  assign llongv[119] = 1'b0;
  assign llongv[118] = 1'b0;
  assign llongv[117] = 1'b0;
  assign llongv[116] = 1'b0;
  assign llongv[115] = 1'b0;
  assign llongv[114] = 1'b0;
  assign llongv[113] = 1'b0;
  assign llongv[112] = 1'b0;
  assign llongv[111] = 1'b0;
  assign llongv[110] = 1'b0;
  assign llongv[109] = 1'b0;
  assign llongv[108] = 1'b0;
  assign llongv[107] = 1'b0;
  assign llongv[106] = 1'b0;
  assign llongv[105] = 1'b0;
  assign llongv[104] = 1'b0;
  assign llongv[103] = 1'b0;
  assign llongv[102] = 1'b0;
  assign llongv[101] = 1'b0;
  assign llongv[100] = 1'b0;
  assign llongv[99] = 1'b0;
  assign llongv[98] = 1'b0;
  assign llongv[97] = 1'b1;
  assign llongv[96] = 1'b0;
  assign llongv[95] = 1'b0;
  assign llongv[94] = 1'b0;
  assign llongv[93] = 1'b0;
  assign llongv[92] = 1'b0;
  assign llongv[91] = 1'b0;
  assign llongv[90] = 1'b0;
  assign llongv[89] = 1'b0;
  assign llongv[88] = 1'b0;
  assign llongv[87] = 1'b0;
  assign llongv[86] = 1'b0;
  assign llongv[85] = 1'b0;
  assign llongv[84] = 1'b0;
  assign llongv[83] = 1'b0;
  assign llongv[82] = 1'b0;
  assign llongv[81] = 1'b0;
  assign llongv[80] = 1'b0;
  assign llongv[79] = 1'b0;
  assign llongv[78] = 1'b0;
  assign llongv[77] = 1'b0;
  assign llongv[76] = 1'b0;
  assign llongv[75] = 1'b0;
  assign llongv[74] = 1'b0;
  assign llongv[73] = 1'b0;
  assign llongv[72] = 1'b0;
  assign llongv[71] = 1'b0;
  assign llongv[70] = 1'b0;
  assign llongv[69] = 1'b0;
  assign llongv[68] = 1'b0;
  assign llongv[67] = 1'b0;
  assign llongv[66] = 1'b0;
  assign llongv[65] = 1'b0;
  assign llongv[64] = 1'b1;
  assign llongv[63] = 1'b0;
  assign llongv[62] = 1'b0;
  assign llongv[61] = 1'b0;
  assign llongv[60] = 1'b0;
  assign llongv[59] = 1'b0;
  assign llongv[58] = 1'b0;
  assign llongv[57] = 1'b0;
  assign llongv[56] = 1'b0;
  assign llongv[55] = 1'b0;
  assign llongv[54] = 1'b0;
  assign llongv[53] = 1'b0;
  assign llongv[52] = 1'b0;
  assign llongv[51] = 1'b0;
  assign llongv[50] = 1'b0;
  assign llongv[49] = 1'b0;
  assign llongv[48] = 1'b0;
  assign llongv[47] = 1'b0;
  assign llongv[46] = 1'b0;
  assign llongv[45] = 1'b0;
  assign llongv[44] = 1'b0;
  assign llongv[43] = 1'b0;
  assign llongv[42] = 1'b0;
  assign llongv[41] = 1'b0;
  assign llongv[40] = 1'b0;
  assign llongv[39] = 1'b0;
  assign llongv[38] = 1'b0;
  assign llongv[37] = 1'b0;
  assign llongv[36] = 1'b0;
  assign llongv[35] = 1'b0;
  assign llongv[34] = 1'b0;
  assign llongv[33] = 1'b1;
  assign llongv[32] = 1'b0;
  assign llongv[31] = 1'b0;
  assign llongv[30] = 1'b0;
  assign llongv[29] = 1'b0;
  assign llongv[28] = 1'b0;
  assign llongv[27] = 1'b0;
  assign llongv[26] = 1'b0;
  assign llongv[25] = 1'b0;
  assign llongv[24] = 1'b0;
  assign llongv[23] = 1'b0;
  assign llongv[22] = 1'b0;
  assign llongv[21] = 1'b0;
  assign llongv[20] = 1'b0;
  assign llongv[19] = 1'b0;
  assign llongv[18] = 1'b0;
  assign llongv[17] = 1'b0;
  assign llongv[16] = 1'b0;
  assign llongv[15] = 1'b0;
  assign llongv[14] = 1'b0;
  assign llongv[13] = 1'b0;
  assign llongv[12] = 1'b0;
  assign llongv[11] = 1'b0;
  assign llongv[10] = 1'b0;
  assign llongv[9] = 1'b0;
  assign llongv[8] = 1'b0;
  assign llongv[7] = 1'b0;
  assign llongv[6] = 1'b0;
  assign llongv[5] = 1'b0;
  assign llongv[4] = 1'b0;
  assign llongv[3] = 1'b0;
  assign llongv[2] = 1'b0;
  assign llongv[1] = 1'b0;
  assign llongv[0] = 1'b1;
  INV_X1_LVT U1_U1_i_0_0 (.ZN(C[0]), .A(A[0]));
  INV_X1_LVT U1_U1_i_0_1 (.ZN(C[1]), .A(B[0]));
  INV_X1_LVT U1_U1_i_0_2 (.ZN(C[2]), .A(B[1]));
  OAI222_X1_LVT U1_U1_i_0_3 (.ZN(C[3]), .A1(A[1]), .A2(A[2]), .B1(B[1]), .B2(
      B[2]), .C1(A[3]), .C2(B[3]));
  INV_X1_LVT U1_U1_i_1_0 (.ZN(C[4]), .A(A[4]));
  INV_X1_LVT U1_U1_i_1_1 (.ZN(C[5]), .A(B[4]));
  INV_X1_LVT U1_U1_i_1_2 (.ZN(C[6]), .A(B[5]));
  OAI222_X1_LVT U1_U1_i_1_3 (.ZN(C[7]), .A1(A[5]), .A2(A[6]), .B1(B[5]), .B2(
      B[6]), .C1(A[7]), .C2(B[7]));
  INV_X1_LVT U1_U1_i_2_0 (.ZN(C[8]), .A(A[8]));
  INV_X1_LVT U1_U1_i_2_1 (.ZN(C[9]), .A(B[8]));
  INV_X1_LVT U1_U1_i_2_2 (.ZN(C[10]), .A(B[9]));
  OAI222_X1_LVT U1_U1_i_2_3 (.ZN(C[11]), .A1(A[9]), .A2(A[10]), .B1(B[9]), .B2(
      B[10]), .C1(A[11]), .C2(B[11]));
  INV_X1_LVT U1_U2_i_0_0 (.ZN(C[12]), .A(A[12]));
  INV_X1_LVT U1_U2_i_0_1 (.ZN(C[13]), .A(B[12]));
  INV_X1_LVT U1_U2_i_0_2 (.ZN(C[14]), .A(B[13]));
  OAI222_X1_LVT U1_U2_i_0_3 (.ZN(C[15]), .A1(A[13]), .A2(A[14]), .B1(B[13]), .B2(
      B[14]), .C1(A[15]), .C2(B[15]));
  INV_X1_LVT U1_U2_i_1_0 (.ZN(C[16]), .A(A[16]));
  INV_X1_LVT U1_U2_i_1_1 (.ZN(C[17]), .A(B[16]));
  INV_X1_LVT U1_U2_i_1_2 (.ZN(C[18]), .A(B[17]));
  OAI222_X1_LVT U1_U2_i_1_3 (.ZN(C[19]), .A1(A[17]), .A2(A[18]), .B1(B[17]), .B2(
      B[18]), .C1(A[19]), .C2(B[19]));
  INV_X1_LVT U1_U2_i_2_0 (.ZN(C[20]), .A(A[20]));
  INV_X1_LVT U1_U2_i_2_1 (.ZN(C[21]), .A(B[20]));
  INV_X1_LVT U1_U2_i_2_2 (.ZN(C[22]), .A(B[21]));
  OAI222_X1_LVT U1_U2_i_2_3 (.ZN(C[23]), .A1(A[21]), .A2(A[22]), .B1(B[21]), .B2(
      B[22]), .C1(A[23]), .C2(B[23]));
  INV_X1_LVT U1_U3_i_0_0 (.ZN(C[24]), .A(A[24]));
  INV_X1_LVT U1_U3_i_0_1 (.ZN(C[25]), .A(B[24]));
  INV_X1_LVT U1_U3_i_0_2 (.ZN(C[26]), .A(B[25]));
  OAI222_X1_LVT U1_U3_i_0_3 (.ZN(C[27]), .A1(A[25]), .A2(A[26]), .B1(B[25]), .B2(
      B[26]), .C1(A[27]), .C2(B[27]));
  INV_X1_LVT U1_U3_i_1_0 (.ZN(C[28]), .A(A[28]));
  INV_X1_LVT U1_U3_i_1_1 (.ZN(C[29]), .A(B[28]));
  INV_X1_LVT U1_U3_i_1_2 (.ZN(C[30]), .A(B[29]));
  OAI222_X1_LVT U1_U3_i_1_3 (.ZN(C[31]), .A1(A[29]), .A2(A[30]), .B1(B[29]), .B2(
      B[30]), .C1(A[31]), .C2(B[31]));
  INV_X1_LVT U1_U3_i_2_0 (.ZN(C[32]), .A(A[32]));
  INV_X1_LVT U1_U3_i_2_1 (.ZN(C[33]), .A(B[32]));
  INV_X1_LVT U1_U3_i_2_2 (.ZN(C[34]), .A(B[33]));
  OAI222_X1_LVT U1_U3_i_2_3 (.ZN(C[35]), .A1(A[33]), .A2(A[34]), .B1(B[33]), .B2(
      B[34]), .C1(A[35]), .C2(B[35]));
  INV_X1_LVT U2_U1_i_0_0 (.ZN(C[41]), .A(A[41]));
  INV_X1_LVT U2_U1_i_0_1 (.ZN(C[42]), .A(B[41]));
  INV_X1_LVT U2_U1_i_0_2 (.ZN(C[43]), .A(B[42]));
  OAI222_X1_LVT U2_U1_i_0_3 (.ZN(C[44]), .A1(A[42]), .A2(A[43]), .B1(B[42]), .B2(
      B[43]), .C1(A[44]), .C2(B[44]));
  INV_X1_LVT U2_U1_i_1_0 (.ZN(C[45]), .A(A[45]));
  INV_X1_LVT U2_U1_i_1_1 (.ZN(C[46]), .A(B[45]));
  INV_X1_LVT U2_U1_i_1_2 (.ZN(C[47]), .A(B[46]));
  OAI222_X1_LVT U2_U1_i_1_3 (.ZN(C[48]), .A1(A[46]), .A2(A[47]), .B1(B[46]), .B2(
      B[47]), .C1(A[48]), .C2(B[48]));
  INV_X1_LVT U2_U1_i_2_0 (.ZN(C[49]), .A(A[49]));
  INV_X1_LVT U2_U1_i_2_1 (.ZN(C[50]), .A(B[49]));
  INV_X1_LVT U2_U1_i_2_2 (.ZN(C[51]), .A(B[50]));
  OAI222_X1_LVT U2_U1_i_2_3 (.ZN(C[52]), .A1(A[50]), .A2(A[51]), .B1(B[50]), .B2(
      B[51]), .C1(A[52]), .C2(B[52]));
  INV_X1_LVT U2_U2_i_0_0 (.ZN(C[53]), .A(A[53]));
  INV_X1_LVT U2_U2_i_0_1 (.ZN(C[54]), .A(B[53]));
  INV_X1_LVT U2_U2_i_0_2 (.ZN(C[55]), .A(B[54]));
  OAI222_X1_LVT U2_U2_i_0_3 (.ZN(C[56]), .A1(A[54]), .A2(A[55]), .B1(B[54]), .B2(
      B[55]), .C1(A[56]), .C2(B[56]));
  INV_X1_LVT U2_U2_i_1_0 (.ZN(C[57]), .A(A[57]));
  INV_X1_LVT U2_U2_i_1_1 (.ZN(C[58]), .A(B[57]));
  INV_X1_LVT U2_U2_i_1_2 (.ZN(C[59]), .A(B[58]));
  OAI222_X1_LVT U2_U2_i_1_3 (.ZN(C[60]), .A1(A[58]), .A2(A[59]), .B1(B[58]), .B2(
      B[59]), .C1(A[60]), .C2(B[60]));
  INV_X1_LVT U2_U2_i_2_0 (.ZN(C[61]), .A(A[61]));
  INV_X1_LVT U2_U2_i_2_1 (.ZN(C[62]), .A(B[61]));
  INV_X1_LVT U2_U2_i_2_2 (.ZN(C[63]), .A(B[62]));
  OAI222_X1_LVT U2_U2_i_2_3 (.ZN(C[64]), .A1(A[62]), .A2(A[63]), .B1(B[62]), .B2(
      B[63]), .C1(A[64]), .C2(B[64]));
  INV_X1_LVT U2_U3_i_0_0 (.ZN(C[65]), .A(A[65]));
  INV_X1_LVT U2_U3_i_0_1 (.ZN(C[66]), .A(B[65]));
  INV_X1_LVT U2_U3_i_0_2 (.ZN(C[67]), .A(B[66]));
  OAI222_X1_LVT U2_U3_i_0_3 (.ZN(C[68]), .A1(A[66]), .A2(A[67]), .B1(B[66]), .B2(
      B[67]), .C1(A[68]), .C2(B[68]));
  INV_X1_LVT U2_U3_i_1_0 (.ZN(C[69]), .A(A[69]));
  INV_X1_LVT U2_U3_i_1_1 (.ZN(C[70]), .A(B[69]));
  INV_X1_LVT U2_U3_i_1_2 (.ZN(C[71]), .A(B[70]));
  OAI222_X1_LVT U2_U3_i_1_3 (.ZN(C[72]), .A1(A[70]), .A2(A[71]), .B1(B[70]), .B2(
      B[71]), .C1(A[72]), .C2(B[72]));
  INV_X1_LVT U2_U3_i_2_0 (.ZN(C[73]), .A(A[73]));
  INV_X1_LVT U2_U3_i_2_1 (.ZN(C[74]), .A(B[73]));
  INV_X1_LVT U2_U3_i_2_2 (.ZN(C[75]), .A(B[74]));
  OAI222_X1_LVT U2_U3_i_2_3 (.ZN(C[76]), .A1(A[74]), .A2(A[75]), .B1(B[74]), .B2(
      B[75]), .C1(A[76]), .C2(B[76]));
  INV_X1_LVT U3_U1_i_0_0 (.ZN(C[82]), .A(1'b1));
  INV_X1_LVT U3_U1_i_0_1 (.ZN(C[83]), .A(longv[41]));
  INV_X1_LVT U3_U1_i_0_2 (.ZN(C[84]), .A(longv[42]));
  OAI222_X1_LVT U3_U1_i_0_3 (.ZN(C[85]), .A1(1'b0), .A2(1'b0), .B1(longv[42]), 
      .B2(longv[43]), .C1(1'b0), .C2(longv[44]));
  INV_X1_LVT U3_U1_i_1_0 (.ZN(C[86]), .A(1'b0));
  INV_X1_LVT U3_U1_i_1_1 (.ZN(C[87]), .A(longv[45]));
  INV_X1_LVT U3_U1_i_1_2 (.ZN(C[88]), .A(longv[46]));
  OAI222_X1_LVT U3_U1_i_1_3 (.ZN(C[89]), .A1(1'b0), .A2(1'b0), .B1(longv[46]), 
      .B2(longv[47]), .C1(1'b0), .C2(longv[48]));
  INV_X1_LVT U3_U1_i_2_0 (.ZN(C[90]), .A(1'b0));
  INV_X1_LVT U3_U1_i_2_1 (.ZN(C[91]), .A(longv[49]));
  INV_X1_LVT U3_U1_i_2_2 (.ZN(C[92]), .A(longv[50]));
  OAI222_X1_LVT U3_U1_i_2_3 (.ZN(C[93]), .A1(1'b0), .A2(1'b0), .B1(longv[50]), 
      .B2(longv[51]), .C1(1'b0), .C2(longv[52]));
  INV_X1_LVT U3_U2_i_0_0 (.ZN(C[94]), .A(1'b0));
  INV_X1_LVT U3_U2_i_0_1 (.ZN(C[95]), .A(longv[53]));
  INV_X1_LVT U3_U2_i_0_2 (.ZN(C[96]), .A(longv[54]));
  OAI222_X1_LVT U3_U2_i_0_3 (.ZN(C[97]), .A1(1'b0), .A2(1'b0), .B1(longv[54]), 
      .B2(longv[55]), .C1(1'b0), .C2(longv[56]));
  INV_X1_LVT U3_U2_i_1_0 (.ZN(C[98]), .A(1'b0));
  INV_X1_LVT U3_U2_i_1_1 (.ZN(C[99]), .A(longv[57]));
  INV_X1_LVT U3_U2_i_1_2 (.ZN(C[100]), .A(longv[58]));
  OAI222_X1_LVT U3_U2_i_1_3 (.ZN(C[101]), .A1(1'b0), .A2(1'b0), .B1(longv[58]), 
      .B2(longv[59]), .C1(1'b0), .C2(longv[60]));
  INV_X1_LVT U3_U2_i_2_0 (.ZN(C[102]), .A(1'b0));
  INV_X1_LVT U3_U2_i_2_1 (.ZN(C[103]), .A(longv[61]));
  INV_X1_LVT U3_U2_i_2_2 (.ZN(C[104]), .A(longv[62]));
  OAI222_X1_LVT U3_U2_i_2_3 (.ZN(C[105]), .A1(1'b0), .A2(1'b0), .B1(longv[62]), 
      .B2(longv[63]), .C1(1'b0), .C2(longv[64]));
  INV_X1_LVT U3_U3_i_0_0 (.ZN(C[106]), .A(1'b0));
  INV_X1_LVT U3_U3_i_0_1 (.ZN(C[107]), .A(longv[65]));
  INV_X1_LVT U3_U3_i_0_2 (.ZN(C[108]), .A(longv[66]));
  OAI222_X1_LVT U3_U3_i_0_3 (.ZN(C[109]), .A1(1'b0), .A2(1'b0), .B1(longv[66]), 
      .B2(longv[67]), .C1(1'b0), .C2(longv[68]));
  INV_X1_LVT U3_U3_i_1_0 (.ZN(C[110]), .A(1'b0));
  INV_X1_LVT U3_U3_i_1_1 (.ZN(C[111]), .A(longv[69]));
  INV_X1_LVT U3_U3_i_1_2 (.ZN(C[112]), .A(longv[70]));
  OAI222_X1_LVT U3_U3_i_1_3 (.ZN(C[113]), .A1(1'b0), .A2(1'b0), .B1(longv[70]), 
      .B2(longv[71]), .C1(1'b0), .C2(longv[72]));
  INV_X1_LVT U3_U3_i_2_0 (.ZN(C[114]), .A(1'b0));
  INV_X1_LVT U3_U3_i_2_1 (.ZN(C[115]), .A(longv[73]));
  INV_X1_LVT U3_U3_i_2_2 (.ZN(C[116]), .A(longv[74]));
  OAI222_X1_LVT U3_U3_i_2_3 (.ZN(C[117]), .A1(1'b1), .A2(1'b0), .B1(longv[74]), 
      .B2(longv[75]), .C1(1'b0), .C2(longv[76]));
endmodule

