module openMSP430(aclk,aclk_en,dbg_freeze,dbg_i2c_sda_out,dbg_uart_txd,
      dco_enable,dco_wkup,dmem_addr,dmem_cen,dmem_din,dmem_wen,irq_acc,
      lfxt_enable,lfxt_wkup,mclk,dma_dout,dma_ready,dma_resp,per_addr,per_din,
      per_en,per_we,pmem_addr,pmem_cen,pmem_din,pmem_wen,puc_rst,smclk,smclk_en,
      cpu_en,dbg_en,dbg_i2c_addr,dbg_i2c_broadcast,dbg_i2c_scl,dbg_i2c_sda_in,
      dbg_uart_rxd,dco_clk,dmem_dout,irq,lfxt_clk,dma_addr,dma_din,dma_en,
      dma_priority,dma_we,dma_wkup,nmi,per_dout,pmem_dout,reset_n,scan_enable,
      scan_mode,wkup);
   output aclk;
   output aclk_en;
   output dbg_freeze;
   output dbg_i2c_sda_out;
   output dbg_uart_txd;
   output dco_enable;
   output dco_wkup;
   output [8:0]dmem_addr;
   output dmem_cen;
   output [15:0]dmem_din;
   output [1:0]dmem_wen;
   output [13:0]irq_acc;
   output lfxt_enable;
   output lfxt_wkup;
   output mclk;
   output [15:0]dma_dout;
   output dma_ready;
   output dma_resp;
   output [13:0]per_addr;
   output [15:0]per_din;
   output per_en;
   output [1:0]per_we;
   output [10:0]pmem_addr;
   output pmem_cen;
   output [15:0]pmem_din;
   output [1:0]pmem_wen;
   output puc_rst;
   output smclk;
   output smclk_en;
   input cpu_en;
   input dbg_en;
   input [6:0]dbg_i2c_addr;
   input [6:0]dbg_i2c_broadcast;
   input dbg_i2c_scl;
   input dbg_i2c_sda_in;
   input dbg_uart_rxd;
   input dco_clk;
   input [15:0]dmem_dout;
   input [13:0]irq;
   input lfxt_clk;
   input [14:0]dma_addr;
   input [15:0]dma_din;
   input dma_en;
   input dma_priority;
   input [1:0]dma_we;
   input dma_wkup;
   input nmi;
   input [15:0]per_dout;
   input [15:0]pmem_dout;
   input reset_n;
   input scan_enable;
   input scan_mode;
   input wkup;
   wire wdtnmies;
   wire wdtifg;
   wire wdt_wkup;
   wire wdt_reset;
   wire wdt_irq;
   wire [15:0]per_dout_wdog;
   wire scg1;
   wire scg0;
   wire pc_sw_wr;
   wire [15:0]pc_sw;
   wire oscoff;
   wire [15:0]eu_mdb_out;
   wire [1:0]eu_mb_wr;
   wire eu_mb_en;
   wire [15:0]eu_mab;
   wire gie;
   wire [15:0]dbg_reg_din;
   wire cpuoff;
   wire [15:0]pc_nxt;
   wire [15:0]pc;
   wire nmi_acc;
   wire mclk_wkup;
   wire mclk_enable;
   wire mclk_dma_wkup;
   wire mclk_dma_enable;
   wire fe_mb_en;
   wire [2:0]inst_type;
   wire [15:0]inst_src;
   wire [7:0]inst_so;
   wire [15:0]inst_sext;
   wire inst_mov;
   wire [7:0]inst_jmp;
   wire inst_irq_rst;
   wire [15:0]inst_dext;
   wire [15:0]inst_dest;
   wire inst_bw;
   wire [11:0]inst_alu;
   wire [7:0]inst_as;
   wire [7:0]inst_ad;
   wire exec_done;
   wire [3:0]e_state;
   wire decode_noirq;
   wire cpu_halt_st;
   wire [15:0]per_dout_mpy;
   wire fe_pmem_wait;
   wire [15:0]fe_mdb_in;
   wire [15:0]eu_mdb_in;
   wire [15:0]dbg_mem_din;
   wire cpu_halt_cmd;
   wire dbg_reg_wr;
   wire [1:0]dbg_mem_wr;
   wire dbg_mem_en;
   wire [15:0]dbg_mem_dout;
   wire [15:0]dbg_mem_addr;
   wire dbg_halt_cmd;
   wire dbg_cpu_reset;
   wire wdtifg_sw_set;
   wire wdtifg_sw_clr;
   wire wdtie;
   wire [15:0]per_dout_sfr;
   wire nmi_wkup;
   wire nmi_pnd;
   wire [31:0]cpu_id;
   wire puc_pnd_set;
   wire por;
   wire [15:0]per_dout_clk;
   wire dbg_rst;
   wire dbg_en_s;
   wire dbg_clk;
   wire cpu_mclk;
   wire cpu_en_s;
   wire n_0_0_0;
   wire [15:0]per_dout_or;
   wire n_0_0_1;
   wire n_0_0_2;
   wire n_0_0_3;
   wire n_0_0_4;
   wire n_0_0_5;
   wire n_0_0_6;
   wire n_0_0_7;
   wire n_0_0_8;
   wire n_0_0_9;
   wire n_0_0_10;
   wire n_0_0_11;
   wire n_0_0_12;
   wire n_0_0_13;
   wire n_0_0_14;
   wire n_0_0_15;
   wire n_14;
   wire n_13;
   wire n_12;
   wire n_11;
   wire n_10;
   wire n_9;
   wire n_8;
   wire n_7;
   wire n_6;
   wire n_5;
   wire n_4;
   wire n_3;
   wire n_2;
   wire n_1;
   wire n_0;
   wire uc_0;
   wire watchdog_0_wdt_rst_noscan;
   wire watchdog_0_wdt_rst;
   wire watchdog_0_wdtcnt_incr;
   wire watchdog_0_wdtcnt_clr_sync;
   wire watchdog_0_wdt_evt_toggle_sync;
   wire watchdog_0_wdt_wkup_pre;
   wire watchdog_0_n_0_0;
   wire watchdog_0_n_0_1;
   wire watchdog_0_n_0_2;
   wire watchdog_0_n_0_3;
   wire watchdog_0_n_0_4;
   wire watchdog_0_reg_wr;
   wire [7:0]watchdog_0_wdtctl;
   wire watchdog_0_n_8_0;
   wire watchdog_0_n_8_1;
   wire watchdog_0_n_8_2;
   wire watchdog_0_wdtpw_error;
   wire watchdog_0_wdt_evt_toggle_sync_dly;
   wire watchdog_0_n_9_0;
   wire watchdog_0_wdtifg_set;
   wire watchdog_0_n_10_0;
   wire watchdog_0_wdtifg_clr;
   wire watchdog_0_n_13_0;
   wire watchdog_0_n_13_1;
   wire watchdog_0_n_17_0;
   wire watchdog_0_wdtcnt_clr_sync_dly;
   wire watchdog_0_n_19_0;
   wire watchdog_0_wdtcnt_clr;
   wire [15:0]watchdog_0_wdtcnt;
   wire watchdog_0_n_21_0;
   wire watchdog_0_n_22_0;
   wire watchdog_0_n_22_1;
   wire [15:0]watchdog_0_wdtcnt_nxt;
   wire watchdog_0_n_24_0;
   wire watchdog_0_n_24_1;
   wire watchdog_0_n_24_2;
   wire watchdog_0_n_24_3;
   wire watchdog_0_n_24_4;
   wire watchdog_0_n_24_5;
   wire watchdog_0_n_24_6;
   wire watchdog_0_n_24_7;
   wire watchdog_0_n_24_8;
   wire watchdog_0_n_24_9;
   wire watchdog_0_n_24_10;
   wire watchdog_0_n_24_11;
   wire watchdog_0_n_24_12;
   wire watchdog_0_n_24_13;
   wire watchdog_0_n_24_14;
   wire [1:0]watchdog_0_wdtisx_ss;
   wire [1:0]watchdog_0_wdtisx_s;
   wire watchdog_0_n_28_0;
   wire watchdog_0_n_28_1;
   wire watchdog_0_n_28_2;
   wire watchdog_0_n_28_3;
   wire watchdog_0_n_28_4;
   wire watchdog_0_n_28_5;
   wire watchdog_0_n_28_6;
   wire watchdog_0_n_28_7;
   wire watchdog_0_n_28_8;
   wire watchdog_0_wdtqn_reg;
   wire watchdog_0_wdtqn_edge;
   wire watchdog_0_wdt_evt_toggle;
   wire watchdog_0_wdt_wkup_en;
   wire watchdog_0_n_35_0;
   wire watchdog_0_n_35_1;
   wire watchdog_0_n_37_0;
   wire watchdog_0_wdtcnt_clr_detect;
   wire watchdog_0_wdtcnt_clr_toggle;
   wire watchdog_0_wdtifg_clr_reg;
   wire watchdog_0_wdtqn_edge_reg;
   wire watchdog_0_n_1;
   wire watchdog_0_n_0;
   wire watchdog_0_n_2;
   wire watchdog_0_n_3;
   wire watchdog_0_n_4;
   wire watchdog_0_n_30;
   wire watchdog_0_n_29;
   wire watchdog_0_n_35;
   wire watchdog_0_n_34;
   wire watchdog_0_n_17;
   wire watchdog_0_n_31;
   wire watchdog_0_n_33;
   wire watchdog_0_n_27;
   wire watchdog_0_n_10;
   wire watchdog_0_n_16;
   wire watchdog_0_n_15;
   wire watchdog_0_n_14;
   wire watchdog_0_n_13;
   wire watchdog_0_n_12;
   wire watchdog_0_n_11;
   wire watchdog_0_n_26;
   wire watchdog_0_n_25;
   wire watchdog_0_n_24;
   wire watchdog_0_n_23;
   wire watchdog_0_n_22;
   wire watchdog_0_n_21;
   wire watchdog_0_n_20;
   wire watchdog_0_n_19;
   wire watchdog_0_n_18;
   wire watchdog_0_n_28;
   wire watchdog_0_n_7;
   wire watchdog_0_n_5;
   wire watchdog_0_n_6;
   wire watchdog_0_n_8;
   wire watchdog_0_n_9;
   wire watchdog_0_n_32;
   wire watchdog_0_sync_reset_por_n_0;
   wire watchdog_0_sync_reset_por_n_1;
   wire watchdog_0_scan_mux_wdt_rst_n_0_0;
   wire watchdog_0_scan_mux_wdt_rst_n_0_1;
   wire watchdog_0_sync_cell_wdtcnt_clr_n_0;
   wire watchdog_0_sync_cell_wdtcnt_clr_n_1;
   wire watchdog_0_sync_cell_wdtcnt_incr_n_0;
   wire watchdog_0_sync_cell_wdtcnt_incr_n_1;
   wire watchdog_0_sync_cell_wdt_evt_n_0;
   wire watchdog_0_sync_cell_wdt_evt_n_1;
   wire watchdog_0_wakeup_cell_wdog_wkup_rst;
   wire watchdog_0_wakeup_cell_wdog_wkup_clk;
   wire watchdog_0_wakeup_cell_wdog_n_0;
   wire watchdog_0_wakeup_cell_wdog_scan_mux_clk_n_0_0;
   wire watchdog_0_wakeup_cell_wdog_scan_mux_clk_n_0_1;
   wire watchdog_0_wakeup_cell_wdog_scan_mux_rst_n_0_0;
   wire watchdog_0_wakeup_cell_wdog_scan_mux_rst_n_0_1;
   wire sfr_0_nmi_capture;
   wire sfr_0_nmi_s;
   wire sfr_0_n_0_0;
   wire sfr_0_n_0_1;
   wire sfr_0_n_0_2;
   wire sfr_0_n_0_3;
   wire sfr_0_reg_sel;
   wire sfr_0_reg_lo_write;
   wire sfr_0_n_2_0;
   wire sfr_0_n_2_1;
   wire sfr_0_n_2_2;
   wire sfr_0_n_2_3;
   wire sfr_0_n_2_4;
   wire sfr_0_n_2_5;
   wire sfr_0_n_2_6;
   wire sfr_0_ifg1_wr;
   wire sfr_0_nmi_capture_rst;
   wire sfr_0_n_4_0;
   wire sfr_0_nmie;
   wire sfr_0_n_7_0;
   wire sfr_0_n_8_0;
   wire sfr_0_n_8_1;
   wire sfr_0_nmi_dly;
   wire sfr_0_n_10_0;
   wire sfr_0_nmi_edge;
   wire sfr_0_nmiifg;
   wire sfr_0_n_13_0;
   wire sfr_0_n_13_1;
   wire sfr_0_n_14_0;
   wire sfr_0_n_14_1;
   wire sfr_0_reg_read;
   wire sfr_0_n_27_0;
   wire sfr_0_n_28_0;
   wire sfr_0_nmi_pol;
   wire sfr_0_n_1;
   wire sfr_0_n_6;
   wire sfr_0_n_11;
   wire sfr_0_n_12;
   wire sfr_0_n_13;
   wire sfr_0_n_10;
   wire sfr_0_n_8;
   wire sfr_0_n_0;
   wire sfr_0_n_5;
   wire sfr_0_n_9;
   wire sfr_0_n_7;
   wire sfr_0_n_31;
   wire sfr_0_n_14;
   wire sfr_0_n_4;
   wire sfr_0_n_19;
   wire sfr_0_n_3;
   wire sfr_0_n_18;
   wire sfr_0_n_25;
   wire sfr_0_n_2;
   wire sfr_0_n_17;
   wire sfr_0_n_24;
   wire sfr_0_n_15;
   wire sfr_0_n_30;
   wire sfr_0_n_16;
   wire sfr_0_n_27;
   wire sfr_0_n_23;
   wire sfr_0_n_22;
   wire sfr_0_n_21;
   wire sfr_0_n_26;
   wire sfr_0_n_20;
   wire sfr_0_n_28;
   wire sfr_0_n_29;
   wire sfr_0_wakeup_cell_nmi_wkup_rst;
   wire sfr_0_wakeup_cell_nmi_wkup_clk;
   wire sfr_0_wakeup_cell_nmi_n_0;
   wire sfr_0_wakeup_cell_nmi_scan_mux_clk_n_0_0;
   wire sfr_0_wakeup_cell_nmi_scan_mux_clk_n_0_1;
   wire sfr_0_wakeup_cell_nmi_scan_mux_rst_n_0_0;
   wire sfr_0_wakeup_cell_nmi_scan_mux_rst_n_0_1;
   wire sfr_0_sync_cell_nmi_n_0;
   wire sfr_0_sync_cell_nmi_n_1;
   wire dbg_0_dbg_wr;
   wire dbg_0_dbg_rd;
   wire [15:0]dbg_0_dbg_din;
   wire [5:0]dbg_0_dbg_addr;
   wire dbg_0_n_0_0;
   wire dbg_0_n_0_1;
   wire dbg_0_n_0_2;
   wire dbg_0_n_0_3;
   wire dbg_0_mem_start;
   wire [2:0]dbg_0_mem_ctl;
   wire dbg_0_mem_burst_rd;
   wire dbg_0_mem_startb;
   wire dbg_0_n_6_0;
   wire dbg_0_n_6_1;
   wire dbg_0_n_8_0;
   wire dbg_0_n_9_0;
   wire dbg_0_n_9_1;
   wire dbg_0_n_9_2;
   wire dbg_0_n_9_3;
   wire dbg_0_n_9_4;
   wire dbg_0_n_9_5;
   wire [1:0]dbg_0_mem_state_nxt_reg;
   wire dbg_0_n_9_6;
   wire [1:0]dbg_0_mem_state;
   wire dbg_0_n_12_0;
   wire dbg_0_mem_access;
   wire dbg_0_n_16_0;
   wire dbg_0_n_17_0;
   wire dbg_0_n_17_1;
   wire dbg_0_n_17_2;
   wire dbg_0_n_17_3;
   wire dbg_0_n_17_4;
   wire dbg_0_n_17_5;
   wire dbg_0_n_17_6;
   wire dbg_0_n_19_0;
   wire dbg_0_n_19_1;
   wire dbg_0_n_19_2;
   wire dbg_0_n_19_3;
   wire dbg_0_n_19_4;
   wire dbg_0_n_19_5;
   wire dbg_0_n_19_6;
   wire dbg_0_n_19_7;
   wire dbg_0_n_19_8;
   wire dbg_0_n_19_9;
   wire dbg_0_n_19_10;
   wire dbg_0_n_19_11;
   wire dbg_0_n_19_12;
   wire dbg_0_n_19_13;
   wire dbg_0_n_19_14;
   wire dbg_0_n_19_15;
   wire dbg_0_n_20_0;
   wire dbg_0_n_20_1;
   wire dbg_0_n_20_2;
   wire dbg_0_n_20_3;
   wire dbg_0_n_20_4;
   wire dbg_0_n_20_5;
   wire dbg_0_n_20_6;
   wire dbg_0_n_20_7;
   wire dbg_0_n_20_8;
   wire dbg_0_n_20_9;
   wire dbg_0_n_20_10;
   wire dbg_0_n_20_11;
   wire dbg_0_n_20_12;
   wire dbg_0_n_20_13;
   wire dbg_0_n_20_14;
   wire dbg_0_n_20_15;
   wire dbg_0_n_20_16;
   wire dbg_0_n_22_0;
   wire dbg_0_dbg_reg_rd;
   wire dbg_0_dbg_mem_rd;
   wire dbg_0_dbg_mem_rd_dly;
   wire dbg_0_dbg_rd_rdy;
   wire dbg_0_n_32_0;
   wire dbg_0_n_32_1;
   wire dbg_0_n_34_0;
   wire dbg_0_dbg_mem_acc;
   wire dbg_0_n_35_0;
   wire dbg_0_n_35_1;
   wire dbg_0_n_37_0;
   wire dbg_0_n_37_1;
   wire dbg_0_n_37_2;
   wire dbg_0_n_37_3;
   wire dbg_0_n_37_4;
   wire [15:0]dbg_0_mem_cnt;
   wire dbg_0_n_39_0;
   wire dbg_0_n_39_1;
   wire dbg_0_n_39_2;
   wire dbg_0_n_39_3;
   wire dbg_0_n_39_4;
   wire dbg_0_n_39_5;
   wire dbg_0_n_39_6;
   wire dbg_0_n_39_7;
   wire dbg_0_n_39_8;
   wire dbg_0_n_39_9;
   wire dbg_0_n_39_10;
   wire dbg_0_n_39_11;
   wire dbg_0_n_39_12;
   wire dbg_0_n_39_13;
   wire dbg_0_n_39_14;
   wire dbg_0_n_39_15;
   wire dbg_0_n_39_16;
   wire dbg_0_n_40_0;
   wire dbg_0_n_40_1;
   wire dbg_0_n_40_2;
   wire dbg_0_n_40_3;
   wire dbg_0_n_40_4;
   wire dbg_0_n_40_5;
   wire dbg_0_n_40_6;
   wire dbg_0_n_40_7;
   wire dbg_0_n_40_8;
   wire dbg_0_n_40_9;
   wire dbg_0_n_40_10;
   wire dbg_0_n_40_11;
   wire dbg_0_n_40_12;
   wire dbg_0_n_40_13;
   wire dbg_0_n_40_14;
   wire dbg_0_n_40_15;
   wire dbg_0_n_40_16;
   wire dbg_0_n_42_0;
   wire dbg_0_n_42_1;
   wire dbg_0_n_42_2;
   wire dbg_0_n_42_3;
   wire dbg_0_mem_burst_start;
   wire dbg_0_n_44_0;
   wire dbg_0_mem_burst_end;
   wire dbg_0_mem_burst;
   wire dbg_0_n_46_0;
   wire dbg_0_n_46_1;
   wire dbg_0_n_48_0;
   wire [5:0]dbg_0_dbg_addr_in;
   wire dbg_0_n_48_1;
   wire dbg_0_n_48_2;
   wire dbg_0_n_49_0;
   wire dbg_0_n_49_1;
   wire dbg_0_n_49_2;
   wire dbg_0_n_49_3;
   wire dbg_0_n_49_4;
   wire dbg_0_n_49_5;
   wire dbg_0_n_49_6;
   wire dbg_0_n_49_7;
   wire dbg_0_n_49_8;
   wire dbg_0_n_49_9;
   wire dbg_0_n_49_10;
   wire dbg_0_n_49_11;
   wire dbg_0_n_49_12;
   wire dbg_0_n_49_13;
   wire dbg_0_n_49_14;
   wire dbg_0_n_49_15;
   wire dbg_0_n_49_16;
   wire dbg_0_n_49_17;
   wire dbg_0_n_49_18;
   wire dbg_0_n_49_19;
   wire dbg_0_n_49_20;
   wire dbg_0_n_49_21;
   wire dbg_0_cpu_ctl_wr;
   wire dbg_0_mem_ctl_wr;
   wire dbg_0_mem_data_wr;
   wire [3:0]dbg_0_cpu_ctl;
   wire dbg_0_n_53_0;
   wire dbg_0_n_53_1;
   wire dbg_0_n_54_0;
   wire dbg_0_n_54_1;
   wire dbg_0_n_54_2;
   wire dbg_0_n_54_3;
   wire dbg_0_n_54_4;
   wire dbg_0_dbg_swbrk;
   wire dbg_0_n_55_0;
   wire dbg_0_n_55_1;
   wire dbg_0_n_55_2;
   wire dbg_0_n_55_3;
   wire dbg_0_n_55_4;
   wire dbg_0_n_55_5;
   wire dbg_0_halt_flag_set;
   wire dbg_0_n_57_0;
   wire dbg_0_n_57_1;
   wire dbg_0_n_57_2;
   wire dbg_0_halt_flag_clr;
   wire dbg_0_halt_flag;
   wire dbg_0_n_59_0;
   wire dbg_0_n_60_0;
   wire dbg_0_n_60_1;
   wire dbg_0_istep;
   wire dbg_0_n_64_0;
   wire dbg_0_n_64_1;
   wire dbg_0_n_66_0;
   wire dbg_0_n_68_0;
   wire dbg_0_n_68_1;
   wire dbg_0_n_68_2;
   wire dbg_0_n_68_3;
   wire dbg_0_n_68_4;
   wire dbg_0_n_68_5;
   wire dbg_0_n_68_6;
   wire dbg_0_n_68_7;
   wire dbg_0_n_68_8;
   wire [15:0]dbg_0_mem_data;
   wire dbg_0_n_70_0;
   wire dbg_0_n_71_0;
   wire dbg_0_n_71_1;
   wire dbg_0_n_71_2;
   wire dbg_0_n_71_3;
   wire dbg_0_n_71_4;
   wire dbg_0_n_71_5;
   wire dbg_0_n_71_6;
   wire dbg_0_n_71_7;
   wire dbg_0_n_71_8;
   wire dbg_0_n_71_9;
   wire dbg_0_n_71_10;
   wire dbg_0_n_71_11;
   wire dbg_0_n_71_12;
   wire dbg_0_n_71_13;
   wire dbg_0_n_71_14;
   wire dbg_0_n_71_15;
   wire dbg_0_n_72_0;
   wire dbg_0_n_72_1;
   wire dbg_0_n_72_2;
   wire dbg_0_n_74_0;
   wire dbg_0_n_74_1;
   wire dbg_0_n_74_2;
   wire dbg_0_n_74_3;
   wire dbg_0_n_74_4;
   wire dbg_0_n_74_5;
   wire dbg_0_n_74_6;
   wire dbg_0_n_74_7;
   wire dbg_0_n_74_8;
   wire dbg_0_n_74_9;
   wire dbg_0_n_74_10;
   wire dbg_0_n_74_11;
   wire dbg_0_n_74_12;
   wire dbg_0_n_74_13;
   wire dbg_0_n_74_14;
   wire dbg_0_n_74_15;
   wire dbg_0_n_74_16;
   wire dbg_0_n_74_17;
   wire dbg_0_n_74_18;
   wire dbg_0_n_74_19;
   wire [1:0]dbg_0_cpu_stat;
   wire dbg_0_n_76_0;
   wire dbg_0_n_76_1;
   wire dbg_0_n_76_2;
   wire dbg_0_n_76_3;
   wire dbg_0_n_76_4;
   wire dbg_0_n_76_5;
   wire dbg_0_n_76_6;
   wire dbg_0_n_78_0;
   wire dbg_0_n_78_1;
   wire dbg_0_n_78_2;
   wire dbg_0_n_78_3;
   wire dbg_0_n_78_4;
   wire dbg_0_n_78_5;
   wire dbg_0_n_78_6;
   wire dbg_0_n_78_7;
   wire [15:0]dbg_0_dbg_dout;
   wire dbg_0_n_78_8;
   wire dbg_0_n_78_9;
   wire dbg_0_n_78_10;
   wire dbg_0_n_78_11;
   wire dbg_0_n_78_12;
   wire dbg_0_n_78_13;
   wire dbg_0_n_78_14;
   wire dbg_0_n_78_15;
   wire dbg_0_n_78_16;
   wire dbg_0_n_78_17;
   wire dbg_0_n_78_18;
   wire dbg_0_n_78_19;
   wire dbg_0_n_78_20;
   wire dbg_0_n_78_21;
   wire dbg_0_n_78_22;
   wire dbg_0_n_78_23;
   wire dbg_0_n_78_24;
   wire dbg_0_n_78_25;
   wire dbg_0_n_78_26;
   wire dbg_0_n_78_27;
   wire dbg_0_n_78_28;
   wire dbg_0_n_78_29;
   wire dbg_0_n_78_30;
   wire dbg_0_n_78_31;
   wire dbg_0_n_78_32;
   wire dbg_0_n_78_33;
   wire dbg_0_n_78_34;
   wire dbg_0_n_78_35;
   wire dbg_0_n_78_36;
   wire dbg_0_n_78_37;
   wire dbg_0_n_78_38;
   wire dbg_0_n_78_39;
   wire dbg_0_n_78_40;
   wire dbg_0_n_78_41;
   wire dbg_0_n_78_42;
   wire dbg_0_n_78_43;
   wire dbg_0_n_78_44;
   wire dbg_0_n_78_45;
   wire dbg_0_n_78_46;
   wire dbg_0_n_78_47;
   wire dbg_0_n_78_48;
   wire dbg_0_n_78_49;
   wire dbg_0_n_78_50;
   wire dbg_0_n_78_51;
   wire dbg_0_n_78_52;
   wire dbg_0_n_78_53;
   wire dbg_0_n_78_54;
   wire dbg_0_n_78_55;
   wire dbg_0_n_78_56;
   wire dbg_0_n_78_57;
   wire dbg_0_n_78_58;
   wire dbg_0_n_78_59;
   wire dbg_0_n_78_60;
   wire dbg_0_n_78_61;
   wire dbg_0_n_78_62;
   wire dbg_0_n_78_63;
   wire dbg_0_n_78_64;
   wire dbg_0_n_78_65;
   wire dbg_0_n_78_66;
   wire dbg_0_n_78_67;
   wire dbg_0_n_78_68;
   wire dbg_0_n_78_69;
   wire dbg_0_n_78_70;
   wire dbg_0_n_78_71;
   wire dbg_0_n_78_72;
   wire dbg_0_n_78_73;
   wire dbg_0_n_78_74;
   wire dbg_0_n_78_75;
   wire dbg_0_n_78_76;
   wire dbg_0_n_78_77;
   wire dbg_0_n_78_78;
   wire dbg_0_n_78_79;
   wire dbg_0_n_78_80;
   wire dbg_0_n_78_81;
   wire dbg_0_n_78_82;
   wire dbg_0_n_78_83;
   wire dbg_0_n_78_84;
   wire dbg_0_n_78_85;
   wire dbg_0_n_78_86;
   wire dbg_0_n_78_87;
   wire dbg_0_n_78_88;
   wire dbg_0_n_78_89;
   wire dbg_0_n_78_90;
   wire dbg_0_n_78_91;
   wire dbg_0_n_78_92;
   wire dbg_0_n_78_93;
   wire dbg_0_n_78_94;
   wire dbg_0_n_78_95;
   wire dbg_0_n_78_96;
   wire dbg_0_n_78_97;
   wire dbg_0_n_78_98;
   wire dbg_0_n_78_99;
   wire dbg_0_n_78_100;
   wire dbg_0_n_78_101;
   wire dbg_0_n_78_102;
   wire dbg_0_n_78_103;
   wire dbg_0_n_78_104;
   wire dbg_0_n_78_105;
   wire dbg_0_n_78_106;
   wire dbg_0_n_78_107;
   wire dbg_0_n_78_108;
   wire dbg_0_n_78_109;
   wire dbg_0_n_78_110;
   wire dbg_0_n_78_111;
   wire dbg_0_n_78_112;
   wire dbg_0_n_78_113;
   wire dbg_0_n_78_114;
   wire dbg_0_n_78_115;
   wire dbg_0_mem_burst_wr;
   wire dbg_0_n_95;
   wire dbg_0_n_1;
   wire dbg_0_n_104;
   wire dbg_0_n_98;
   wire dbg_0_n_102;
   wire dbg_0_n_55;
   wire dbg_0_n_57;
   wire dbg_0_n_73;
   wire dbg_0_n_58;
   wire dbg_0_n_74;
   wire dbg_0_n_59;
   wire dbg_0_n_75;
   wire dbg_0_n_60;
   wire dbg_0_n_76;
   wire dbg_0_n_61;
   wire dbg_0_n_77;
   wire dbg_0_n_62;
   wire dbg_0_n_78;
   wire dbg_0_n_63;
   wire dbg_0_n_79;
   wire dbg_0_n_64;
   wire dbg_0_n_80;
   wire dbg_0_n_65;
   wire dbg_0_n_81;
   wire dbg_0_n_66;
   wire dbg_0_n_82;
   wire dbg_0_n_67;
   wire dbg_0_n_83;
   wire dbg_0_n_68;
   wire dbg_0_n_84;
   wire dbg_0_n_69;
   wire dbg_0_n_85;
   wire dbg_0_n_70;
   wire dbg_0_n_86;
   wire dbg_0_n_71;
   wire dbg_0_n_87;
   wire dbg_0_n_2;
   wire dbg_0_n_3;
   wire dbg_0_n_4;
   wire dbg_0_n_0;
   wire dbg_0_n_5;
   wire dbg_0_n_6;
   wire dbg_0_n_7;
   wire dbg_0_n_47;
   wire dbg_0_n_48;
   wire dbg_0_n_96;
   wire dbg_0_n_101;
   wire dbg_0_n_10;
   wire dbg_0_n_53;
   wire dbg_0_n_11;
   wire dbg_0_n_13;
   wire dbg_0_n_29;
   wire dbg_0_n_46;
   wire dbg_0_n_45;
   wire dbg_0_n_49;
   wire dbg_0_n_51;
   wire dbg_0_n_9;
   wire dbg_0_n_50;
   wire dbg_0_n_52;
   wire dbg_0_n_54;
   wire dbg_0_n_56;
   wire dbg_0_n_72;
   wire dbg_0_n_88;
   wire dbg_0_n_90;
   wire dbg_0_n_89;
   wire dbg_0_n_27;
   wire dbg_0_n_43;
   wire dbg_0_n_26;
   wire dbg_0_n_42;
   wire dbg_0_n_25;
   wire dbg_0_n_41;
   wire dbg_0_n_24;
   wire dbg_0_n_40;
   wire dbg_0_n_23;
   wire dbg_0_n_39;
   wire dbg_0_n_22;
   wire dbg_0_n_38;
   wire dbg_0_n_21;
   wire dbg_0_n_37;
   wire dbg_0_n_20;
   wire dbg_0_n_36;
   wire dbg_0_n_19;
   wire dbg_0_n_35;
   wire dbg_0_n_18;
   wire dbg_0_n_34;
   wire dbg_0_n_17;
   wire dbg_0_n_33;
   wire dbg_0_n_16;
   wire dbg_0_n_32;
   wire dbg_0_n_15;
   wire dbg_0_n_31;
   wire dbg_0_n_12;
   wire dbg_0_n_14;
   wire dbg_0_n_30;
   wire dbg_0_n_28;
   wire dbg_0_n_44;
   wire dbg_0_n_97;
   wire dbg_0_n_136;
   wire dbg_0_n_135;
   wire dbg_0_n_115;
   wire dbg_0_n_133;
   wire dbg_0_n_152;
   wire dbg_0_n_153;
   wire dbg_0_n_134;
   wire dbg_0_n_92;
   wire dbg_0_n_91;
   wire dbg_0_n_99;
   wire dbg_0_n_132;
   wire dbg_0_n_151;
   wire dbg_0_n_131;
   wire dbg_0_n_150;
   wire dbg_0_n_130;
   wire dbg_0_n_149;
   wire dbg_0_n_129;
   wire dbg_0_n_148;
   wire dbg_0_n_128;
   wire dbg_0_n_147;
   wire dbg_0_n_127;
   wire dbg_0_n_146;
   wire dbg_0_n_126;
   wire dbg_0_n_145;
   wire dbg_0_n_116;
   wire dbg_0_n_117;
   wire dbg_0_n_125;
   wire dbg_0_n_144;
   wire dbg_0_n_124;
   wire dbg_0_n_143;
   wire dbg_0_n_93;
   wire dbg_0_n_123;
   wire dbg_0_n_142;
   wire dbg_0_n_105;
   wire dbg_0_n_122;
   wire dbg_0_n_141;
   wire dbg_0_n_106;
   wire dbg_0_n_121;
   wire dbg_0_n_140;
   wire dbg_0_n_94;
   wire dbg_0_n_107;
   wire dbg_0_n_100;
   wire dbg_0_n_155;
   wire dbg_0_n_120;
   wire dbg_0_n_139;
   wire dbg_0_n_154;
   wire dbg_0_n_119;
   wire dbg_0_n_138;
   wire dbg_0_n_118;
   wire dbg_0_n_137;
   wire dbg_0_n_103;
   wire dbg_0_n_8;
   wire dbg_0_n_108;
   wire dbg_0_n_110;
   wire dbg_0_n_111;
   wire dbg_0_n_109;
   wire dbg_0_n_113;
   wire dbg_0_n_114;
   wire dbg_0_n_112;
   wire dbg_0_dbg_uart_0_uart_rxd_n;
   wire dbg_0_dbg_uart_0_uart_rxd;
   wire [1:0]dbg_0_dbg_uart_0_rxd_buf;
   wire dbg_0_dbg_uart_0_n_2_0;
   wire dbg_0_dbg_uart_0_n_2_1;
   wire dbg_0_dbg_uart_0_n_2_2;
   wire dbg_0_dbg_uart_0_rxd_maj_nxt;
   wire [19:0]dbg_0_dbg_uart_0_xfer_buf;
   wire dbg_0_dbg_uart_0_n_4_0;
   wire dbg_0_dbg_uart_0_n_4_1;
   wire dbg_0_dbg_uart_0_n_4_2;
   wire dbg_0_dbg_uart_0_n_4_3;
   wire dbg_0_dbg_uart_0_n_4_4;
   wire dbg_0_dbg_uart_0_n_4_5;
   wire dbg_0_dbg_uart_0_n_4_6;
   wire dbg_0_dbg_uart_0_n_4_7;
   wire dbg_0_dbg_uart_0_n_4_8;
   wire dbg_0_dbg_uart_0_n_4_9;
   wire dbg_0_dbg_uart_0_n_4_10;
   wire dbg_0_dbg_uart_0_n_4_11;
   wire dbg_0_dbg_uart_0_n_4_12;
   wire dbg_0_dbg_uart_0_n_4_13;
   wire dbg_0_dbg_uart_0_n_4_14;
   wire dbg_0_dbg_uart_0_n_4_15;
   wire dbg_0_dbg_uart_0_n_4_16;
   wire dbg_0_dbg_uart_0_n_4_17;
   wire dbg_0_dbg_uart_0_n_4_18;
   wire dbg_0_dbg_uart_0_n_5_0;
   wire dbg_0_dbg_uart_0_n_5_1;
   wire dbg_0_dbg_uart_0_rxd_maj;
   wire dbg_0_dbg_uart_0_n_7_0;
   wire dbg_0_dbg_uart_0_n_8_0;
   wire dbg_0_dbg_uart_0_n_8_1;
   wire dbg_0_dbg_uart_0_n_8_2;
   wire dbg_0_dbg_uart_0_n_8_3;
   wire dbg_0_dbg_uart_0_n_8_4;
   wire dbg_0_dbg_uart_0_n_8_5;
   wire dbg_0_dbg_uart_0_n_8_6;
   wire dbg_0_dbg_uart_0_n_8_7;
   wire dbg_0_dbg_uart_0_n_8_8;
   wire dbg_0_dbg_uart_0_n_8_9;
   wire dbg_0_dbg_uart_0_n_8_10;
   wire dbg_0_dbg_uart_0_n_8_11;
   wire dbg_0_dbg_uart_0_n_8_12;
   wire dbg_0_dbg_uart_0_n_8_13;
   wire dbg_0_dbg_uart_0_n_8_14;
   wire dbg_0_dbg_uart_0_n_8_15;
   wire dbg_0_dbg_uart_0_n_8_16;
   wire dbg_0_dbg_uart_0_n_8_17;
   wire dbg_0_dbg_uart_0_n_8_18;
   wire dbg_0_dbg_uart_0_n_8_19;
   wire dbg_0_dbg_uart_0_n_8_20;
   wire dbg_0_dbg_uart_0_n_8_21;
   wire dbg_0_dbg_uart_0_n_8_22;
   wire dbg_0_dbg_uart_0_n_8_23;
   wire dbg_0_dbg_uart_0_n_8_24;
   wire [2:0]dbg_0_dbg_uart_0_uart_state_nxt_reg;
   wire dbg_0_dbg_uart_0_n_8_25;
   wire dbg_0_dbg_uart_0_n_8_26;
   wire dbg_0_dbg_uart_0_n_8_27;
   wire dbg_0_dbg_uart_0_n_8_28;
   wire dbg_0_dbg_uart_0_n_8_29;
   wire [2:0]dbg_0_dbg_uart_0_uart_state;
   wire dbg_0_dbg_uart_0_n_11_0;
   wire dbg_0_dbg_uart_0_n_11_1;
   wire dbg_0_dbg_uart_0_n_13_0;
   wire dbg_0_dbg_uart_0_n_13_1;
   wire dbg_0_dbg_uart_0_n_13_2;
   wire dbg_0_dbg_uart_0_n_14_0;
   wire dbg_0_dbg_uart_0_n_15_0;
   wire dbg_0_dbg_uart_0_rxd_fe;
   wire dbg_0_dbg_uart_0_sync_busy;
   wire [15:0]dbg_0_dbg_uart_0_bit_cnt_max;
   wire dbg_0_dbg_uart_0_n_21_0;
   wire dbg_0_dbg_uart_0_n_21_1;
   wire dbg_0_dbg_uart_0_n_21_2;
   wire dbg_0_dbg_uart_0_n_21_3;
   wire dbg_0_dbg_uart_0_n_21_4;
   wire dbg_0_dbg_uart_0_n_21_5;
   wire dbg_0_dbg_uart_0_n_21_6;
   wire dbg_0_dbg_uart_0_n_21_7;
   wire dbg_0_dbg_uart_0_n_21_8;
   wire dbg_0_dbg_uart_0_n_21_9;
   wire dbg_0_dbg_uart_0_n_21_10;
   wire dbg_0_dbg_uart_0_n_21_11;
   wire dbg_0_dbg_uart_0_n_21_12;
   wire dbg_0_dbg_uart_0_n_21_13;
   wire dbg_0_dbg_uart_0_n_21_14;
   wire dbg_0_dbg_uart_0_n_21_15;
   wire dbg_0_dbg_uart_0_n_21_16;
   wire dbg_0_dbg_uart_0_n_21_17;
   wire dbg_0_dbg_uart_0_n_22_0;
   wire dbg_0_dbg_uart_0_n_22_1;
   wire dbg_0_dbg_uart_0_n_24_0;
   wire dbg_0_dbg_uart_0_txd_start;
   wire dbg_0_dbg_uart_0_rx_active;
   wire [15:0]dbg_0_dbg_uart_0_xfer_cnt;
   wire dbg_0_dbg_uart_0_n_27_0;
   wire dbg_0_dbg_uart_0_n_27_1;
   wire dbg_0_dbg_uart_0_n_27_2;
   wire dbg_0_dbg_uart_0_n_27_3;
   wire dbg_0_dbg_uart_0_n_27_4;
   wire dbg_0_dbg_uart_0_n_27_5;
   wire dbg_0_dbg_uart_0_n_27_6;
   wire dbg_0_dbg_uart_0_n_27_7;
   wire dbg_0_dbg_uart_0_n_27_8;
   wire dbg_0_dbg_uart_0_n_27_9;
   wire dbg_0_dbg_uart_0_n_27_10;
   wire dbg_0_dbg_uart_0_n_27_11;
   wire dbg_0_dbg_uart_0_n_27_12;
   wire dbg_0_dbg_uart_0_n_27_13;
   wire dbg_0_dbg_uart_0_n_29_0;
   wire dbg_0_dbg_uart_0_n_30_0;
   wire dbg_0_dbg_uart_0_n_31_0;
   wire dbg_0_dbg_uart_0_n_31_1;
   wire dbg_0_dbg_uart_0_n_31_2;
   wire dbg_0_dbg_uart_0_n_31_3;
   wire dbg_0_dbg_uart_0_n_31_4;
   wire dbg_0_dbg_uart_0_n_31_5;
   wire dbg_0_dbg_uart_0_n_31_6;
   wire dbg_0_dbg_uart_0_n_31_7;
   wire dbg_0_dbg_uart_0_n_31_8;
   wire dbg_0_dbg_uart_0_n_31_9;
   wire dbg_0_dbg_uart_0_n_31_10;
   wire dbg_0_dbg_uart_0_n_31_11;
   wire dbg_0_dbg_uart_0_n_31_12;
   wire dbg_0_dbg_uart_0_n_31_13;
   wire dbg_0_dbg_uart_0_n_31_14;
   wire dbg_0_dbg_uart_0_n_31_15;
   wire dbg_0_dbg_uart_0_n_31_16;
   wire dbg_0_dbg_uart_0_n_31_17;
   wire dbg_0_dbg_uart_0_n_31_18;
   wire dbg_0_dbg_uart_0_n_31_19;
   wire dbg_0_dbg_uart_0_n_31_20;
   wire dbg_0_dbg_uart_0_n_31_21;
   wire dbg_0_dbg_uart_0_n_31_22;
   wire dbg_0_dbg_uart_0_n_31_23;
   wire dbg_0_dbg_uart_0_n_31_24;
   wire dbg_0_dbg_uart_0_n_31_25;
   wire dbg_0_dbg_uart_0_n_31_26;
   wire dbg_0_dbg_uart_0_n_31_27;
   wire dbg_0_dbg_uart_0_n_31_28;
   wire dbg_0_dbg_uart_0_n_31_29;
   wire dbg_0_dbg_uart_0_n_31_30;
   wire dbg_0_dbg_uart_0_n_31_31;
   wire dbg_0_dbg_uart_0_n_31_32;
   wire dbg_0_dbg_uart_0_n_32_0;
   wire dbg_0_dbg_uart_0_n_32_1;
   wire dbg_0_dbg_uart_0_n_32_2;
   wire dbg_0_dbg_uart_0_n_32_3;
   wire dbg_0_dbg_uart_0_n_33_0;
   wire dbg_0_dbg_uart_0_n_33_1;
   wire dbg_0_dbg_uart_0_n_33_2;
   wire dbg_0_dbg_uart_0_n_35_0;
   wire dbg_0_dbg_uart_0_n_35_1;
   wire dbg_0_dbg_uart_0_n_35_2;
   wire dbg_0_dbg_uart_0_n_35_3;
   wire dbg_0_dbg_uart_0_n_35_4;
   wire dbg_0_dbg_uart_0_n_35_5;
   wire dbg_0_dbg_uart_0_xfer_bit_inc;
   wire [3:0]dbg_0_dbg_uart_0_xfer_bit;
   wire dbg_0_dbg_uart_0_n_39_0;
   wire dbg_0_dbg_uart_0_n_39_1;
   wire dbg_0_dbg_uart_0_n_39_2;
   wire dbg_0_dbg_uart_0_n_40_0;
   wire dbg_0_dbg_uart_0_n_41_0;
   wire dbg_0_dbg_uart_0_n_41_1;
   wire dbg_0_dbg_uart_0_n_42_0;
   wire dbg_0_dbg_uart_0_n_42_1;
   wire dbg_0_dbg_uart_0_n_42_2;
   wire dbg_0_dbg_uart_0_n_44_0;
   wire dbg_0_dbg_uart_0_n_44_1;
   wire dbg_0_dbg_uart_0_n_44_2;
   wire dbg_0_dbg_uart_0_n_44_3;
   wire dbg_0_dbg_uart_0_xfer_done;
   wire dbg_0_dbg_uart_0_cmd_valid;
   wire dbg_0_dbg_uart_0_dbg_bw;
   wire dbg_0_dbg_uart_0_n_49_0;
   wire dbg_0_dbg_uart_0_n_49_1;
   wire dbg_0_dbg_uart_0_n_49_2;
   wire dbg_0_dbg_uart_0_n_49_3;
   wire dbg_0_dbg_uart_0_n_49_4;
   wire dbg_0_dbg_uart_0_n_49_5;
   wire dbg_0_dbg_uart_0_n_49_6;
   wire dbg_0_dbg_uart_0_n_49_7;
   wire dbg_0_dbg_uart_0_n_49_8;
   wire dbg_0_dbg_uart_0_n_49_9;
   wire dbg_0_dbg_uart_0_n_49_10;
   wire dbg_0_dbg_uart_0_n_50_0;
   wire dbg_0_dbg_uart_0_n_50_1;
   wire dbg_0_dbg_uart_0_n_52_0;
   wire dbg_0_dbg_uart_0_n_52_1;
   wire dbg_0_dbg_uart_0_n_54_0;
   wire dbg_0_dbg_uart_0_n_136;
   wire dbg_0_dbg_uart_0_n_130;
   wire dbg_0_dbg_uart_0_n_19;
   wire dbg_0_dbg_uart_0_n_76;
   wire dbg_0_dbg_uart_0_n_53;
   wire dbg_0_dbg_uart_0_n_58;
   wire dbg_0_dbg_uart_0_n_54;
   wire dbg_0_dbg_uart_0_n_56;
   wire dbg_0_dbg_uart_0_n_57;
   wire dbg_0_dbg_uart_0_n_55;
   wire dbg_0_dbg_uart_0_n_52;
   wire dbg_0_dbg_uart_0_n_59;
   wire dbg_0_dbg_uart_0_n_51;
   wire dbg_0_dbg_uart_0_n_22;
   wire dbg_0_dbg_uart_0_n_119;
   wire dbg_0_dbg_uart_0_n_123;
   wire dbg_0_dbg_uart_0_n_124;
   wire dbg_0_dbg_uart_0_n_128;
   wire dbg_0_dbg_uart_0_n_118;
   wire dbg_0_dbg_uart_0_n_120;
   wire dbg_0_dbg_uart_0_n_125;
   wire dbg_0_dbg_uart_0_n_121;
   wire dbg_0_dbg_uart_0_n_122;
   wire dbg_0_dbg_uart_0_n_127;
   wire dbg_0_dbg_uart_0_n_116;
   wire dbg_0_dbg_uart_0_n_117;
   wire dbg_0_dbg_uart_0_n_28;
   wire dbg_0_dbg_uart_0_n_126;
   wire dbg_0_dbg_uart_0_n_25;
   wire dbg_0_dbg_uart_0_n_27;
   wire dbg_0_dbg_uart_0_n_26;
   wire dbg_0_dbg_uart_0_n_29;
   wire dbg_0_dbg_uart_0_n_31;
   wire dbg_0_dbg_uart_0_n_24;
   wire dbg_0_dbg_uart_0_n_23;
   wire dbg_0_dbg_uart_0_n_33;
   wire dbg_0_dbg_uart_0_n_34;
   wire dbg_0_dbg_uart_0_n_32;
   wire dbg_0_dbg_uart_0_n_50;
   wire dbg_0_dbg_uart_0_n_60;
   wire dbg_0_dbg_uart_0_n_61;
   wire dbg_0_dbg_uart_0_n_49;
   wire dbg_0_dbg_uart_0_n_95;
   wire dbg_0_dbg_uart_0_n_94;
   wire dbg_0_dbg_uart_0_n_97;
   wire dbg_0_dbg_uart_0_n_78;
   wire dbg_0_dbg_uart_0_n_96;
   wire dbg_0_dbg_uart_0_n_98;
   wire dbg_0_dbg_uart_0_n_79;
   wire dbg_0_dbg_uart_0_n_62;
   wire dbg_0_dbg_uart_0_n_48;
   wire dbg_0_dbg_uart_0_n_99;
   wire dbg_0_dbg_uart_0_n_77;
   wire dbg_0_dbg_uart_0_n_80;
   wire dbg_0_dbg_uart_0_n_63;
   wire dbg_0_dbg_uart_0_n_47;
   wire dbg_0_dbg_uart_0_n_100;
   wire dbg_0_dbg_uart_0_n_81;
   wire dbg_0_dbg_uart_0_n_64;
   wire dbg_0_dbg_uart_0_n_46;
   wire dbg_0_dbg_uart_0_n_101;
   wire dbg_0_dbg_uart_0_n_82;
   wire dbg_0_dbg_uart_0_n_65;
   wire dbg_0_dbg_uart_0_n_45;
   wire dbg_0_dbg_uart_0_n_102;
   wire dbg_0_dbg_uart_0_n_83;
   wire dbg_0_dbg_uart_0_n_66;
   wire dbg_0_dbg_uart_0_n_44;
   wire dbg_0_dbg_uart_0_n_103;
   wire dbg_0_dbg_uart_0_n_84;
   wire dbg_0_dbg_uart_0_n_67;
   wire dbg_0_dbg_uart_0_n_43;
   wire dbg_0_dbg_uart_0_n_104;
   wire dbg_0_dbg_uart_0_n_85;
   wire dbg_0_dbg_uart_0_n_68;
   wire dbg_0_dbg_uart_0_n_42;
   wire dbg_0_dbg_uart_0_n_105;
   wire dbg_0_dbg_uart_0_n_86;
   wire dbg_0_dbg_uart_0_n_69;
   wire dbg_0_dbg_uart_0_n_41;
   wire dbg_0_dbg_uart_0_n_106;
   wire dbg_0_dbg_uart_0_n_87;
   wire dbg_0_dbg_uart_0_n_70;
   wire dbg_0_dbg_uart_0_n_40;
   wire dbg_0_dbg_uart_0_n_107;
   wire dbg_0_dbg_uart_0_n_88;
   wire dbg_0_dbg_uart_0_n_71;
   wire dbg_0_dbg_uart_0_n_39;
   wire dbg_0_dbg_uart_0_n_108;
   wire dbg_0_dbg_uart_0_n_89;
   wire dbg_0_dbg_uart_0_n_72;
   wire dbg_0_dbg_uart_0_n_38;
   wire dbg_0_dbg_uart_0_n_109;
   wire dbg_0_dbg_uart_0_n_90;
   wire dbg_0_dbg_uart_0_n_73;
   wire dbg_0_dbg_uart_0_n_37;
   wire dbg_0_dbg_uart_0_n_110;
   wire dbg_0_dbg_uart_0_n_91;
   wire dbg_0_dbg_uart_0_n_74;
   wire dbg_0_dbg_uart_0_n_36;
   wire dbg_0_dbg_uart_0_n_111;
   wire dbg_0_dbg_uart_0_n_92;
   wire dbg_0_dbg_uart_0_n_75;
   wire dbg_0_dbg_uart_0_n_35;
   wire dbg_0_dbg_uart_0_n_112;
   wire dbg_0_dbg_uart_0_n_93;
   wire dbg_0_dbg_uart_0_n_113;
   wire dbg_0_dbg_uart_0_n_114;
   wire dbg_0_dbg_uart_0_n_115;
   wire dbg_0_dbg_uart_0_n_21;
   wire dbg_0_dbg_uart_0_n_0;
   wire dbg_0_dbg_uart_0_n_18;
   wire dbg_0_dbg_uart_0_n_17;
   wire dbg_0_dbg_uart_0_n_129;
   wire dbg_0_dbg_uart_0_n_16;
   wire dbg_0_dbg_uart_0_n_15;
   wire dbg_0_dbg_uart_0_n_14;
   wire dbg_0_dbg_uart_0_n_13;
   wire dbg_0_dbg_uart_0_n_12;
   wire dbg_0_dbg_uart_0_n_131;
   wire dbg_0_dbg_uart_0_n_11;
   wire dbg_0_dbg_uart_0_n_10;
   wire dbg_0_dbg_uart_0_n_20;
   wire dbg_0_dbg_uart_0_n_9;
   wire dbg_0_dbg_uart_0_n_8;
   wire dbg_0_dbg_uart_0_n_7;
   wire dbg_0_dbg_uart_0_n_6;
   wire dbg_0_dbg_uart_0_n_5;
   wire dbg_0_dbg_uart_0_n_4;
   wire dbg_0_dbg_uart_0_n_132;
   wire dbg_0_dbg_uart_0_n_30;
   wire dbg_0_dbg_uart_0_n_133;
   wire dbg_0_dbg_uart_0_n_3;
   wire dbg_0_dbg_uart_0_n_2;
   wire dbg_0_dbg_uart_0_n_1;
   wire dbg_0_dbg_uart_0_n_135;
   wire dbg_0_dbg_uart_0_n_134;
   wire dbg_0_dbg_uart_0_sync_cell_uart_rxd_n_0;
   wire dbg_0_dbg_uart_0_sync_cell_uart_rxd_n_1;
   wire multiplier_0_n_0_0;
   wire multiplier_0_n_0_1;
   wire multiplier_0_n_0_2;
   wire multiplier_0_n_0_3;
   wire multiplier_0_reg_sel;
   wire multiplier_0_reg_read;
   wire multiplier_0_n_3_0;
   wire multiplier_0_n_3_1;
   wire multiplier_0_n_3_2;
   wire multiplier_0_reg_rd1;
   wire multiplier_0_reg_rd15;
   wire multiplier_0_reg_write;
   wire multiplier_0_op2_wr;
   wire multiplier_0_reslo_wr;
   wire multiplier_0_reshi_wr;
   wire [15:0]multiplier_0_per_din_msk;
   wire [15:0]multiplier_0_op2_reg;
   wire [1:0]multiplier_0_cycle;
   wire multiplier_0_result_wr;
   wire multiplier_0_op1_wr;
   wire multiplier_0_sign_sel;
   wire [8:0]multiplier_0_op2_hi_xp;
   wire multiplier_0_n_29_0;
   wire multiplier_0_n_29_1;
   wire [8:0]multiplier_0_op2_xp;
   wire multiplier_0_n_29_2;
   wire multiplier_0_n_29_3;
   wire multiplier_0_n_29_4;
   wire multiplier_0_n_29_5;
   wire multiplier_0_n_29_6;
   wire multiplier_0_n_29_7;
   wire multiplier_0_n_29_8;
   wire [15:0]multiplier_0_op1;
   wire [16:0]multiplier_0_op1_xp;
   wire multiplier_0_n_32_0;
   wire multiplier_0_n_32_1;
   wire multiplier_0_n_32_2;
   wire multiplier_0_n_32_3;
   wire multiplier_0_n_32_4;
   wire multiplier_0_n_32_5;
   wire multiplier_0_n_32_6;
   wire multiplier_0_n_32_7;
   wire multiplier_0_n_32_8;
   wire multiplier_0_n_32_9;
   wire multiplier_0_n_32_10;
   wire multiplier_0_n_32_11;
   wire multiplier_0_n_32_12;
   wire multiplier_0_n_32_13;
   wire multiplier_0_n_32_14;
   wire multiplier_0_n_32_15;
   wire multiplier_0_n_32_16;
   wire multiplier_0_n_32_17;
   wire multiplier_0_n_32_18;
   wire multiplier_0_n_32_19;
   wire multiplier_0_n_32_20;
   wire multiplier_0_n_32_21;
   wire multiplier_0_n_32_22;
   wire multiplier_0_n_32_23;
   wire multiplier_0_n_32_24;
   wire multiplier_0_n_32_25;
   wire multiplier_0_n_32_26;
   wire multiplier_0_n_32_27;
   wire multiplier_0_n_32_28;
   wire multiplier_0_n_32_29;
   wire multiplier_0_n_32_30;
   wire multiplier_0_n_32_31;
   wire multiplier_0_n_32_32;
   wire multiplier_0_n_32_33;
   wire multiplier_0_n_32_34;
   wire multiplier_0_n_32_35;
   wire multiplier_0_n_32_36;
   wire multiplier_0_n_32_37;
   wire multiplier_0_n_32_38;
   wire multiplier_0_n_32_39;
   wire multiplier_0_n_32_40;
   wire multiplier_0_n_32_41;
   wire multiplier_0_n_32_42;
   wire multiplier_0_n_32_43;
   wire multiplier_0_n_32_44;
   wire multiplier_0_n_32_45;
   wire multiplier_0_n_32_46;
   wire multiplier_0_n_32_47;
   wire multiplier_0_n_32_48;
   wire multiplier_0_n_32_49;
   wire multiplier_0_n_32_50;
   wire multiplier_0_n_32_51;
   wire multiplier_0_n_32_52;
   wire multiplier_0_n_32_53;
   wire multiplier_0_n_32_54;
   wire multiplier_0_n_32_55;
   wire multiplier_0_n_32_56;
   wire multiplier_0_n_32_57;
   wire multiplier_0_n_32_58;
   wire multiplier_0_n_32_59;
   wire multiplier_0_n_32_60;
   wire multiplier_0_n_32_61;
   wire multiplier_0_n_32_62;
   wire multiplier_0_n_32_63;
   wire multiplier_0_n_32_64;
   wire multiplier_0_n_32_65;
   wire multiplier_0_n_32_66;
   wire multiplier_0_n_32_67;
   wire multiplier_0_n_32_68;
   wire multiplier_0_n_32_69;
   wire multiplier_0_n_32_70;
   wire multiplier_0_n_32_71;
   wire multiplier_0_n_32_72;
   wire multiplier_0_n_32_73;
   wire multiplier_0_n_32_74;
   wire multiplier_0_n_32_75;
   wire multiplier_0_n_32_76;
   wire multiplier_0_n_32_77;
   wire multiplier_0_n_32_78;
   wire multiplier_0_n_32_79;
   wire multiplier_0_n_32_80;
   wire multiplier_0_n_32_81;
   wire multiplier_0_n_32_82;
   wire multiplier_0_n_32_83;
   wire multiplier_0_n_32_84;
   wire multiplier_0_n_32_85;
   wire multiplier_0_n_32_86;
   wire multiplier_0_n_32_87;
   wire multiplier_0_n_32_88;
   wire multiplier_0_n_32_89;
   wire multiplier_0_n_32_90;
   wire multiplier_0_n_32_91;
   wire multiplier_0_n_32_92;
   wire multiplier_0_n_32_93;
   wire multiplier_0_n_32_94;
   wire multiplier_0_n_32_95;
   wire multiplier_0_n_32_96;
   wire multiplier_0_n_32_97;
   wire multiplier_0_n_32_98;
   wire multiplier_0_n_32_99;
   wire multiplier_0_n_32_100;
   wire multiplier_0_n_32_101;
   wire multiplier_0_n_32_102;
   wire multiplier_0_n_32_103;
   wire multiplier_0_n_32_104;
   wire multiplier_0_n_32_105;
   wire multiplier_0_n_32_106;
   wire multiplier_0_n_32_107;
   wire multiplier_0_n_32_108;
   wire multiplier_0_n_32_109;
   wire multiplier_0_n_32_110;
   wire multiplier_0_n_32_111;
   wire multiplier_0_n_32_112;
   wire multiplier_0_n_32_113;
   wire multiplier_0_n_32_114;
   wire multiplier_0_n_32_115;
   wire multiplier_0_n_32_116;
   wire multiplier_0_n_32_117;
   wire multiplier_0_n_32_118;
   wire multiplier_0_n_32_119;
   wire multiplier_0_n_32_120;
   wire multiplier_0_n_32_121;
   wire multiplier_0_n_32_122;
   wire multiplier_0_n_32_123;
   wire multiplier_0_n_32_124;
   wire multiplier_0_n_32_125;
   wire multiplier_0_n_32_126;
   wire multiplier_0_n_32_127;
   wire multiplier_0_n_32_128;
   wire multiplier_0_n_32_129;
   wire multiplier_0_n_32_130;
   wire multiplier_0_n_32_131;
   wire multiplier_0_n_32_132;
   wire multiplier_0_n_32_133;
   wire multiplier_0_n_32_134;
   wire multiplier_0_n_32_135;
   wire multiplier_0_n_32_136;
   wire multiplier_0_n_32_137;
   wire multiplier_0_n_32_138;
   wire multiplier_0_n_32_139;
   wire multiplier_0_n_32_140;
   wire multiplier_0_n_32_141;
   wire multiplier_0_n_32_142;
   wire multiplier_0_n_32_143;
   wire multiplier_0_n_32_144;
   wire multiplier_0_n_32_145;
   wire multiplier_0_n_32_146;
   wire multiplier_0_n_32_147;
   wire multiplier_0_n_32_148;
   wire multiplier_0_n_32_149;
   wire multiplier_0_n_32_150;
   wire multiplier_0_n_32_151;
   wire multiplier_0_n_32_152;
   wire multiplier_0_n_32_153;
   wire multiplier_0_n_32_154;
   wire multiplier_0_n_32_155;
   wire multiplier_0_n_32_156;
   wire multiplier_0_n_32_157;
   wire multiplier_0_n_32_158;
   wire multiplier_0_n_32_159;
   wire multiplier_0_n_32_160;
   wire multiplier_0_n_32_161;
   wire multiplier_0_n_32_162;
   wire multiplier_0_n_32_163;
   wire multiplier_0_n_32_164;
   wire multiplier_0_n_32_165;
   wire multiplier_0_n_32_166;
   wire multiplier_0_n_32_167;
   wire multiplier_0_n_32_168;
   wire multiplier_0_n_32_169;
   wire multiplier_0_n_32_170;
   wire multiplier_0_n_32_171;
   wire multiplier_0_n_32_172;
   wire multiplier_0_n_32_173;
   wire multiplier_0_n_32_174;
   wire multiplier_0_n_32_175;
   wire multiplier_0_n_32_176;
   wire multiplier_0_n_32_177;
   wire multiplier_0_n_32_178;
   wire multiplier_0_n_32_179;
   wire multiplier_0_n_32_180;
   wire multiplier_0_n_32_181;
   wire multiplier_0_n_32_182;
   wire multiplier_0_n_32_183;
   wire multiplier_0_n_32_184;
   wire multiplier_0_n_32_185;
   wire multiplier_0_n_32_186;
   wire multiplier_0_n_32_187;
   wire multiplier_0_n_32_188;
   wire multiplier_0_n_32_189;
   wire multiplier_0_n_32_190;
   wire multiplier_0_n_32_191;
   wire multiplier_0_n_32_192;
   wire multiplier_0_n_32_193;
   wire multiplier_0_n_32_194;
   wire multiplier_0_n_32_195;
   wire multiplier_0_n_32_196;
   wire multiplier_0_n_32_197;
   wire multiplier_0_n_32_198;
   wire multiplier_0_n_32_199;
   wire multiplier_0_n_32_200;
   wire multiplier_0_n_32_201;
   wire multiplier_0_n_32_202;
   wire multiplier_0_n_32_203;
   wire multiplier_0_n_32_204;
   wire multiplier_0_n_32_205;
   wire multiplier_0_n_32_206;
   wire multiplier_0_n_32_207;
   wire multiplier_0_n_32_208;
   wire multiplier_0_n_32_209;
   wire multiplier_0_n_32_210;
   wire multiplier_0_n_32_211;
   wire multiplier_0_n_32_212;
   wire multiplier_0_n_32_213;
   wire multiplier_0_n_32_214;
   wire multiplier_0_n_32_215;
   wire multiplier_0_n_32_216;
   wire multiplier_0_n_32_217;
   wire multiplier_0_n_32_218;
   wire multiplier_0_n_32_219;
   wire multiplier_0_n_32_220;
   wire multiplier_0_n_32_221;
   wire multiplier_0_n_32_222;
   wire multiplier_0_n_32_223;
   wire multiplier_0_n_32_224;
   wire multiplier_0_n_32_225;
   wire multiplier_0_n_32_226;
   wire multiplier_0_n_32_227;
   wire multiplier_0_n_32_228;
   wire multiplier_0_n_32_229;
   wire multiplier_0_n_32_230;
   wire multiplier_0_n_32_231;
   wire multiplier_0_n_32_232;
   wire multiplier_0_n_32_233;
   wire multiplier_0_n_32_234;
   wire multiplier_0_n_32_235;
   wire multiplier_0_n_32_236;
   wire multiplier_0_n_32_237;
   wire multiplier_0_n_32_238;
   wire multiplier_0_n_32_239;
   wire multiplier_0_n_32_240;
   wire multiplier_0_n_32_241;
   wire multiplier_0_n_32_242;
   wire multiplier_0_n_32_243;
   wire multiplier_0_n_32_244;
   wire multiplier_0_n_32_245;
   wire multiplier_0_n_32_246;
   wire multiplier_0_n_32_247;
   wire multiplier_0_n_32_248;
   wire multiplier_0_n_32_249;
   wire multiplier_0_n_32_250;
   wire multiplier_0_n_32_251;
   wire multiplier_0_n_32_252;
   wire multiplier_0_n_32_253;
   wire multiplier_0_n_32_254;
   wire multiplier_0_n_32_255;
   wire multiplier_0_n_32_256;
   wire multiplier_0_n_32_257;
   wire multiplier_0_n_32_258;
   wire multiplier_0_n_32_259;
   wire multiplier_0_n_32_260;
   wire multiplier_0_n_32_261;
   wire multiplier_0_n_32_262;
   wire multiplier_0_n_32_263;
   wire multiplier_0_n_32_264;
   wire multiplier_0_n_32_265;
   wire multiplier_0_n_32_266;
   wire multiplier_0_n_32_267;
   wire multiplier_0_n_32_268;
   wire multiplier_0_n_32_269;
   wire multiplier_0_n_32_270;
   wire multiplier_0_n_32_271;
   wire multiplier_0_n_32_272;
   wire multiplier_0_n_32_273;
   wire multiplier_0_n_32_274;
   wire multiplier_0_n_32_275;
   wire multiplier_0_n_32_276;
   wire multiplier_0_n_32_277;
   wire multiplier_0_n_32_278;
   wire multiplier_0_n_32_279;
   wire multiplier_0_n_32_280;
   wire multiplier_0_n_32_281;
   wire multiplier_0_n_32_282;
   wire multiplier_0_n_32_283;
   wire multiplier_0_n_32_284;
   wire multiplier_0_n_32_285;
   wire multiplier_0_n_32_286;
   wire multiplier_0_n_32_287;
   wire multiplier_0_n_32_288;
   wire multiplier_0_n_32_289;
   wire multiplier_0_n_32_290;
   wire multiplier_0_n_32_291;
   wire multiplier_0_n_32_292;
   wire multiplier_0_n_32_293;
   wire multiplier_0_n_32_294;
   wire multiplier_0_n_32_295;
   wire multiplier_0_n_32_296;
   wire multiplier_0_n_32_297;
   wire multiplier_0_n_32_298;
   wire multiplier_0_n_32_299;
   wire multiplier_0_n_32_300;
   wire multiplier_0_n_32_301;
   wire multiplier_0_n_32_302;
   wire multiplier_0_n_32_303;
   wire multiplier_0_n_32_304;
   wire multiplier_0_n_32_305;
   wire multiplier_0_n_32_306;
   wire multiplier_0_n_32_307;
   wire multiplier_0_n_32_308;
   wire multiplier_0_n_32_309;
   wire multiplier_0_n_32_310;
   wire multiplier_0_n_32_311;
   wire multiplier_0_n_32_312;
   wire multiplier_0_n_32_313;
   wire multiplier_0_n_32_314;
   wire multiplier_0_n_32_315;
   wire multiplier_0_n_32_316;
   wire multiplier_0_n_32_317;
   wire multiplier_0_n_32_318;
   wire multiplier_0_n_32_319;
   wire multiplier_0_n_32_320;
   wire multiplier_0_n_32_321;
   wire multiplier_0_n_32_322;
   wire multiplier_0_n_32_323;
   wire multiplier_0_n_32_324;
   wire multiplier_0_n_32_325;
   wire multiplier_0_n_32_326;
   wire multiplier_0_n_32_327;
   wire multiplier_0_n_32_328;
   wire multiplier_0_n_32_329;
   wire multiplier_0_n_32_330;
   wire multiplier_0_n_32_331;
   wire multiplier_0_n_32_332;
   wire multiplier_0_n_32_333;
   wire multiplier_0_n_32_334;
   wire multiplier_0_n_32_335;
   wire multiplier_0_n_32_336;
   wire multiplier_0_n_32_337;
   wire multiplier_0_n_32_338;
   wire multiplier_0_n_32_339;
   wire multiplier_0_n_32_340;
   wire multiplier_0_n_32_341;
   wire multiplier_0_n_32_342;
   wire multiplier_0_n_32_343;
   wire multiplier_0_n_32_344;
   wire multiplier_0_n_32_345;
   wire multiplier_0_n_32_346;
   wire multiplier_0_n_32_347;
   wire multiplier_0_n_32_348;
   wire multiplier_0_n_32_349;
   wire multiplier_0_n_32_350;
   wire multiplier_0_n_32_351;
   wire multiplier_0_n_32_352;
   wire multiplier_0_n_32_353;
   wire multiplier_0_n_32_354;
   wire multiplier_0_n_32_355;
   wire multiplier_0_n_32_356;
   wire multiplier_0_n_32_357;
   wire multiplier_0_n_32_358;
   wire multiplier_0_n_32_359;
   wire multiplier_0_n_32_360;
   wire multiplier_0_n_32_361;
   wire multiplier_0_n_32_362;
   wire multiplier_0_n_32_363;
   wire multiplier_0_n_32_364;
   wire multiplier_0_n_32_365;
   wire multiplier_0_n_32_366;
   wire multiplier_0_n_32_367;
   wire multiplier_0_n_32_368;
   wire multiplier_0_n_32_369;
   wire multiplier_0_n_32_370;
   wire multiplier_0_n_32_371;
   wire multiplier_0_n_32_372;
   wire multiplier_0_n_32_373;
   wire multiplier_0_n_32_374;
   wire multiplier_0_n_32_375;
   wire multiplier_0_n_32_376;
   wire multiplier_0_n_32_377;
   wire multiplier_0_n_32_378;
   wire multiplier_0_n_32_379;
   wire multiplier_0_n_32_380;
   wire multiplier_0_n_32_381;
   wire multiplier_0_n_32_382;
   wire multiplier_0_n_32_383;
   wire multiplier_0_n_32_384;
   wire multiplier_0_n_32_385;
   wire multiplier_0_n_32_386;
   wire multiplier_0_n_32_387;
   wire multiplier_0_n_32_388;
   wire multiplier_0_n_32_389;
   wire multiplier_0_n_32_390;
   wire multiplier_0_n_32_391;
   wire multiplier_0_n_32_392;
   wire multiplier_0_n_32_393;
   wire multiplier_0_n_32_394;
   wire multiplier_0_n_32_395;
   wire multiplier_0_n_32_396;
   wire multiplier_0_n_32_397;
   wire multiplier_0_n_32_398;
   wire multiplier_0_n_32_399;
   wire multiplier_0_n_32_400;
   wire multiplier_0_n_32_401;
   wire multiplier_0_n_32_402;
   wire multiplier_0_n_32_403;
   wire multiplier_0_n_32_404;
   wire multiplier_0_n_32_405;
   wire multiplier_0_n_32_406;
   wire multiplier_0_n_32_407;
   wire multiplier_0_n_32_408;
   wire multiplier_0_n_32_409;
   wire multiplier_0_n_32_410;
   wire multiplier_0_n_32_411;
   wire multiplier_0_n_32_412;
   wire multiplier_0_n_32_413;
   wire multiplier_0_n_32_414;
   wire multiplier_0_n_32_415;
   wire multiplier_0_n_32_416;
   wire multiplier_0_n_32_417;
   wire multiplier_0_n_32_418;
   wire multiplier_0_n_32_419;
   wire multiplier_0_n_32_420;
   wire multiplier_0_n_32_421;
   wire multiplier_0_n_32_422;
   wire multiplier_0_n_32_423;
   wire multiplier_0_n_32_424;
   wire multiplier_0_n_32_425;
   wire multiplier_0_n_32_426;
   wire multiplier_0_n_32_427;
   wire multiplier_0_n_32_428;
   wire multiplier_0_n_32_429;
   wire multiplier_0_n_32_430;
   wire multiplier_0_n_32_431;
   wire multiplier_0_n_32_432;
   wire multiplier_0_n_32_433;
   wire multiplier_0_n_32_434;
   wire multiplier_0_n_32_435;
   wire multiplier_0_n_32_436;
   wire multiplier_0_n_32_437;
   wire multiplier_0_n_32_438;
   wire multiplier_0_n_32_439;
   wire multiplier_0_n_32_440;
   wire multiplier_0_n_32_441;
   wire multiplier_0_n_32_442;
   wire multiplier_0_n_32_443;
   wire multiplier_0_n_32_444;
   wire multiplier_0_n_32_445;
   wire multiplier_0_n_32_446;
   wire multiplier_0_n_32_447;
   wire multiplier_0_n_32_448;
   wire multiplier_0_n_32_449;
   wire multiplier_0_n_32_450;
   wire multiplier_0_n_32_451;
   wire multiplier_0_n_32_452;
   wire multiplier_0_n_32_453;
   wire multiplier_0_n_32_454;
   wire multiplier_0_n_32_455;
   wire multiplier_0_n_32_456;
   wire multiplier_0_n_32_457;
   wire multiplier_0_n_32_458;
   wire multiplier_0_n_32_459;
   wire multiplier_0_n_32_460;
   wire multiplier_0_n_32_461;
   wire multiplier_0_n_32_462;
   wire multiplier_0_n_32_463;
   wire multiplier_0_n_32_464;
   wire multiplier_0_n_32_465;
   wire multiplier_0_n_32_466;
   wire multiplier_0_n_32_467;
   wire multiplier_0_n_32_468;
   wire multiplier_0_n_32_469;
   wire multiplier_0_n_32_470;
   wire multiplier_0_n_32_471;
   wire multiplier_0_n_32_472;
   wire multiplier_0_n_32_473;
   wire multiplier_0_n_32_474;
   wire multiplier_0_n_32_475;
   wire multiplier_0_n_32_476;
   wire multiplier_0_n_32_477;
   wire multiplier_0_n_32_478;
   wire multiplier_0_n_32_479;
   wire multiplier_0_n_32_480;
   wire multiplier_0_n_32_481;
   wire multiplier_0_n_32_482;
   wire multiplier_0_n_32_483;
   wire multiplier_0_n_32_484;
   wire multiplier_0_n_32_485;
   wire multiplier_0_n_32_486;
   wire multiplier_0_n_32_487;
   wire multiplier_0_n_32_488;
   wire multiplier_0_n_32_489;
   wire multiplier_0_n_32_490;
   wire multiplier_0_n_32_491;
   wire multiplier_0_n_32_492;
   wire multiplier_0_n_32_493;
   wire multiplier_0_n_32_494;
   wire multiplier_0_n_32_495;
   wire multiplier_0_n_32_496;
   wire multiplier_0_n_32_497;
   wire multiplier_0_n_32_498;
   wire multiplier_0_n_32_499;
   wire multiplier_0_n_32_500;
   wire multiplier_0_n_32_501;
   wire multiplier_0_n_32_502;
   wire multiplier_0_n_32_503;
   wire multiplier_0_n_32_504;
   wire multiplier_0_n_32_505;
   wire multiplier_0_n_32_506;
   wire multiplier_0_n_32_507;
   wire multiplier_0_n_32_508;
   wire multiplier_0_n_32_509;
   wire multiplier_0_n_32_510;
   wire multiplier_0_n_32_511;
   wire multiplier_0_n_32_512;
   wire multiplier_0_n_32_513;
   wire multiplier_0_n_32_514;
   wire multiplier_0_n_32_515;
   wire multiplier_0_n_32_516;
   wire multiplier_0_n_32_517;
   wire multiplier_0_n_32_518;
   wire multiplier_0_n_32_519;
   wire multiplier_0_n_32_520;
   wire multiplier_0_n_32_521;
   wire multiplier_0_n_32_522;
   wire multiplier_0_n_32_523;
   wire multiplier_0_n_32_524;
   wire multiplier_0_n_32_525;
   wire multiplier_0_n_32_526;
   wire multiplier_0_n_32_527;
   wire multiplier_0_n_32_528;
   wire multiplier_0_n_32_529;
   wire multiplier_0_n_32_530;
   wire multiplier_0_n_32_531;
   wire multiplier_0_n_32_532;
   wire multiplier_0_n_32_533;
   wire multiplier_0_n_32_534;
   wire multiplier_0_n_32_535;
   wire multiplier_0_n_32_536;
   wire multiplier_0_n_32_537;
   wire multiplier_0_n_32_538;
   wire multiplier_0_n_32_539;
   wire multiplier_0_n_32_540;
   wire multiplier_0_n_32_541;
   wire multiplier_0_n_32_542;
   wire multiplier_0_n_32_543;
   wire multiplier_0_n_32_544;
   wire multiplier_0_n_32_545;
   wire multiplier_0_n_32_546;
   wire multiplier_0_n_32_547;
   wire multiplier_0_n_32_548;
   wire multiplier_0_n_32_549;
   wire multiplier_0_n_32_550;
   wire multiplier_0_n_32_551;
   wire multiplier_0_n_32_552;
   wire multiplier_0_n_32_553;
   wire multiplier_0_n_32_554;
   wire multiplier_0_n_32_555;
   wire multiplier_0_n_32_556;
   wire multiplier_0_n_32_557;
   wire multiplier_0_n_32_558;
   wire multiplier_0_n_32_559;
   wire multiplier_0_n_32_560;
   wire multiplier_0_n_32_561;
   wire multiplier_0_n_32_562;
   wire multiplier_0_n_32_563;
   wire multiplier_0_n_32_564;
   wire multiplier_0_n_32_565;
   wire multiplier_0_n_32_566;
   wire multiplier_0_n_32_567;
   wire multiplier_0_n_32_568;
   wire multiplier_0_n_32_569;
   wire multiplier_0_n_32_570;
   wire multiplier_0_n_32_571;
   wire multiplier_0_n_32_572;
   wire multiplier_0_n_32_573;
   wire multiplier_0_n_32_574;
   wire multiplier_0_n_32_575;
   wire multiplier_0_n_32_576;
   wire multiplier_0_n_32_577;
   wire multiplier_0_n_32_578;
   wire multiplier_0_n_32_579;
   wire multiplier_0_n_32_580;
   wire multiplier_0_n_32_581;
   wire multiplier_0_n_32_582;
   wire multiplier_0_n_32_583;
   wire multiplier_0_n_32_584;
   wire multiplier_0_n_32_585;
   wire multiplier_0_n_32_586;
   wire multiplier_0_n_32_587;
   wire multiplier_0_n_32_588;
   wire multiplier_0_n_32_589;
   wire multiplier_0_n_32_590;
   wire multiplier_0_n_32_591;
   wire multiplier_0_n_32_592;
   wire multiplier_0_n_32_593;
   wire multiplier_0_n_32_594;
   wire multiplier_0_n_32_595;
   wire multiplier_0_n_32_596;
   wire multiplier_0_n_32_597;
   wire multiplier_0_n_32_598;
   wire multiplier_0_n_32_599;
   wire multiplier_0_n_32_600;
   wire multiplier_0_n_32_601;
   wire multiplier_0_n_32_602;
   wire multiplier_0_n_32_603;
   wire multiplier_0_n_32_604;
   wire multiplier_0_n_32_605;
   wire multiplier_0_n_32_606;
   wire multiplier_0_n_32_607;
   wire multiplier_0_n_32_608;
   wire multiplier_0_n_32_609;
   wire multiplier_0_n_32_610;
   wire multiplier_0_n_32_611;
   wire multiplier_0_n_32_612;
   wire multiplier_0_n_32_613;
   wire multiplier_0_n_32_614;
   wire multiplier_0_n_32_615;
   wire multiplier_0_n_32_616;
   wire multiplier_0_n_32_617;
   wire multiplier_0_n_32_618;
   wire multiplier_0_n_32_619;
   wire multiplier_0_n_32_620;
   wire multiplier_0_n_32_621;
   wire multiplier_0_n_32_622;
   wire multiplier_0_n_32_623;
   wire multiplier_0_n_32_624;
   wire multiplier_0_n_32_625;
   wire multiplier_0_n_32_626;
   wire multiplier_0_n_32_627;
   wire multiplier_0_n_32_628;
   wire multiplier_0_n_32_629;
   wire multiplier_0_n_32_630;
   wire multiplier_0_n_32_631;
   wire multiplier_0_n_32_632;
   wire multiplier_0_n_32_633;
   wire multiplier_0_n_32_634;
   wire multiplier_0_n_32_635;
   wire multiplier_0_n_32_636;
   wire multiplier_0_n_32_637;
   wire multiplier_0_n_32_638;
   wire multiplier_0_n_32_639;
   wire multiplier_0_n_32_640;
   wire multiplier_0_n_32_641;
   wire multiplier_0_n_32_642;
   wire multiplier_0_n_32_643;
   wire multiplier_0_n_32_644;
   wire multiplier_0_n_32_645;
   wire multiplier_0_n_32_646;
   wire multiplier_0_n_32_647;
   wire multiplier_0_n_32_648;
   wire multiplier_0_n_32_649;
   wire multiplier_0_n_32_650;
   wire multiplier_0_n_32_651;
   wire multiplier_0_n_32_652;
   wire multiplier_0_n_32_653;
   wire multiplier_0_n_32_654;
   wire multiplier_0_n_32_655;
   wire multiplier_0_n_32_656;
   wire multiplier_0_n_32_657;
   wire multiplier_0_n_32_658;
   wire multiplier_0_n_32_659;
   wire multiplier_0_n_32_660;
   wire multiplier_0_n_32_661;
   wire multiplier_0_n_32_662;
   wire multiplier_0_n_32_663;
   wire multiplier_0_n_32_664;
   wire multiplier_0_n_32_665;
   wire multiplier_0_n_32_666;
   wire multiplier_0_n_32_667;
   wire multiplier_0_n_32_668;
   wire multiplier_0_n_32_669;
   wire multiplier_0_n_32_670;
   wire multiplier_0_n_32_671;
   wire multiplier_0_n_32_672;
   wire multiplier_0_n_32_673;
   wire multiplier_0_n_32_674;
   wire multiplier_0_n_34_0;
   wire [31:0]multiplier_0_product_xp;
   wire multiplier_0_n_34_1;
   wire multiplier_0_n_34_2;
   wire multiplier_0_n_34_3;
   wire multiplier_0_n_34_4;
   wire multiplier_0_n_34_5;
   wire multiplier_0_n_34_6;
   wire multiplier_0_n_34_7;
   wire multiplier_0_n_34_8;
   wire multiplier_0_n_34_9;
   wire multiplier_0_n_34_10;
   wire multiplier_0_n_34_11;
   wire multiplier_0_n_34_12;
   wire multiplier_0_n_34_13;
   wire multiplier_0_n_34_14;
   wire multiplier_0_n_34_15;
   wire multiplier_0_n_34_16;
   wire multiplier_0_n_34_17;
   wire multiplier_0_n_34_18;
   wire multiplier_0_n_34_19;
   wire multiplier_0_n_34_20;
   wire multiplier_0_n_34_21;
   wire multiplier_0_n_34_22;
   wire multiplier_0_n_34_23;
   wire multiplier_0_n_34_24;
   wire multiplier_0_n_34_25;
   wire multiplier_0_acc_sel;
   wire multiplier_0_n_38_0;
   wire multiplier_0_result_clr;
   wire multiplier_0_n_39_0;
   wire multiplier_0_n_39_1;
   wire [15:0]multiplier_0_reshi;
   wire multiplier_0_n_41_0;
   wire multiplier_0_n_41_1;
   wire multiplier_0_n_41_2;
   wire multiplier_0_n_41_3;
   wire multiplier_0_n_41_4;
   wire multiplier_0_n_41_5;
   wire multiplier_0_n_41_6;
   wire multiplier_0_n_41_7;
   wire multiplier_0_n_41_8;
   wire multiplier_0_n_41_9;
   wire multiplier_0_n_41_10;
   wire multiplier_0_n_41_11;
   wire multiplier_0_n_41_12;
   wire multiplier_0_n_41_13;
   wire multiplier_0_n_41_14;
   wire multiplier_0_n_41_15;
   wire multiplier_0_n_41_16;
   wire multiplier_0_n_42_0;
   wire multiplier_0_n_42_1;
   wire multiplier_0_n_45_0;
   wire multiplier_0_n_45_1;
   wire multiplier_0_n_45_2;
   wire multiplier_0_n_45_3;
   wire multiplier_0_n_45_4;
   wire multiplier_0_n_45_5;
   wire multiplier_0_n_45_6;
   wire multiplier_0_n_45_7;
   wire multiplier_0_n_45_8;
   wire multiplier_0_n_45_9;
   wire multiplier_0_n_45_10;
   wire multiplier_0_n_45_11;
   wire multiplier_0_n_45_12;
   wire multiplier_0_n_45_13;
   wire multiplier_0_n_45_14;
   wire multiplier_0_n_45_15;
   wire multiplier_0_n_45_16;
   wire multiplier_0_n_46_0;
   wire multiplier_0_n_46_1;
   wire multiplier_0_n_48_0;
   wire multiplier_0_n_48_1;
   wire multiplier_0_n_48_2;
   wire multiplier_0_n_48_3;
   wire multiplier_0_n_48_4;
   wire multiplier_0_n_48_5;
   wire multiplier_0_n_48_6;
   wire multiplier_0_n_48_7;
   wire multiplier_0_n_48_8;
   wire multiplier_0_n_48_9;
   wire multiplier_0_n_48_10;
   wire multiplier_0_n_48_11;
   wire multiplier_0_n_48_12;
   wire multiplier_0_n_48_13;
   wire multiplier_0_n_48_14;
   wire multiplier_0_n_48_15;
   wire [15:0]multiplier_0_reshi_nxt;
   wire multiplier_0_n_48_16;
   wire multiplier_0_n_48_17;
   wire multiplier_0_n_48_18;
   wire multiplier_0_n_48_19;
   wire multiplier_0_n_48_20;
   wire multiplier_0_n_48_21;
   wire multiplier_0_n_48_22;
   wire multiplier_0_n_48_23;
   wire multiplier_0_n_48_24;
   wire multiplier_0_n_48_25;
   wire multiplier_0_n_48_26;
   wire multiplier_0_n_48_27;
   wire multiplier_0_n_48_28;
   wire multiplier_0_n_48_29;
   wire multiplier_0_n_48_30;
   wire multiplier_0_n_50_0;
   wire multiplier_0_n_50_1;
   wire [1:0]multiplier_0_sumext_s_nxt;
   wire [1:0]multiplier_0_sumext_s;
   wire multiplier_0_n_52_0;
   wire multiplier_0_n_53_0;
   wire multiplier_0_n_53_1;
   wire multiplier_0_n_55_0;
   wire multiplier_0_n_55_1;
   wire multiplier_0_n_55_2;
   wire multiplier_0_n_57_0;
   wire multiplier_0_n_57_1;
   wire multiplier_0_n_60_0;
   wire multiplier_0_n_60_1;
   wire multiplier_0_n_60_2;
   wire multiplier_0_n_60_3;
   wire multiplier_0_n_60_4;
   wire multiplier_0_n_60_5;
   wire multiplier_0_n_60_6;
   wire multiplier_0_n_60_7;
   wire multiplier_0_n_60_8;
   wire multiplier_0_n_60_9;
   wire multiplier_0_n_60_10;
   wire multiplier_0_n_60_11;
   wire multiplier_0_n_60_12;
   wire multiplier_0_n_60_13;
   wire multiplier_0_n_60_14;
   wire multiplier_0_n_60_15;
   wire multiplier_0_n_60_16;
   wire multiplier_0_n_60_17;
   wire multiplier_0_n_60_18;
   wire multiplier_0_n_60_19;
   wire multiplier_0_n_60_20;
   wire multiplier_0_n_60_21;
   wire multiplier_0_n_60_22;
   wire multiplier_0_n_60_23;
   wire multiplier_0_n_60_24;
   wire multiplier_0_n_60_25;
   wire multiplier_0_n_60_26;
   wire multiplier_0_n_60_27;
   wire multiplier_0_n_60_28;
   wire multiplier_0_n_60_29;
   wire multiplier_0_n_60_30;
   wire multiplier_0_n_60_31;
   wire multiplier_0_n_60_32;
   wire multiplier_0_n_60_33;
   wire multiplier_0_n_60_34;
   wire multiplier_0_n_60_35;
   wire multiplier_0_n_60_36;
   wire multiplier_0_n_60_37;
   wire multiplier_0_n_60_38;
   wire multiplier_0_n_60_39;
   wire multiplier_0_n_60_40;
   wire multiplier_0_n_60_41;
   wire multiplier_0_n_60_42;
   wire multiplier_0_n_60_43;
   wire multiplier_0_n_60_44;
   wire multiplier_0_n_60_45;
   wire multiplier_0_n_60_46;
   wire multiplier_0_n_60_47;
   wire multiplier_0_n_60_48;
   wire multiplier_0_n_60_49;
   wire multiplier_0_n_60_50;
   wire multiplier_0_n_60_51;
   wire multiplier_0_n_60_52;
   wire multiplier_0_n_60_53;
   wire multiplier_0_n_60_54;
   wire multiplier_0_n_60_55;
   wire multiplier_0_n_60_56;
   wire multiplier_0_n_60_57;
   wire multiplier_0_n_60_58;
   wire multiplier_0_n_60_59;
   wire multiplier_0_n_60_60;
   wire multiplier_0_n_60_61;
   wire multiplier_0_n_60_62;
   wire multiplier_0_n_60_63;
   wire multiplier_0_n_60_64;
   wire multiplier_0_n_60_65;
   wire multiplier_0_n_60_66;
   wire multiplier_0_n_60_67;
   wire multiplier_0_n_60_68;
   wire multiplier_0_n_60_69;
   wire multiplier_0_n_60_70;
   wire multiplier_0_n_60_71;
   wire multiplier_0_n_60_72;
   wire multiplier_0_n_60_73;
   wire multiplier_0_n_60_74;
   wire multiplier_0_n_60_75;
   wire multiplier_0_n_60_76;
   wire multiplier_0_n_60_77;
   wire multiplier_0_n_60_78;
   wire multiplier_0_n_60_79;
   wire multiplier_0_n_60_80;
   wire multiplier_0_n_60_81;
   wire multiplier_0_n_60_82;
   wire multiplier_0_n_15;
   wire multiplier_0_n_5;
   wire multiplier_0_n_38;
   wire multiplier_0_n_3;
   wire multiplier_0_n_18;
   wire multiplier_0_n_4;
   wire multiplier_0_n_19;
   wire multiplier_0_n_68;
   wire multiplier_0_n_1;
   wire multiplier_0_n_16;
   wire multiplier_0_n_2;
   wire multiplier_0_n_17;
   wire multiplier_0_n_67;
   wire multiplier_0_n_6;
   wire multiplier_0_n_20;
   wire multiplier_0_n_21;
   wire multiplier_0_n_41;
   wire multiplier_0_n_45;
   wire multiplier_0_n_46;
   wire multiplier_0_n_47;
   wire multiplier_0_n_48;
   wire multiplier_0_n_49;
   wire multiplier_0_n_40;
   wire multiplier_0_n_39;
   wire multiplier_0_n_50;
   wire multiplier_0_n_51;
   wire multiplier_0_n_52;
   wire multiplier_0_n_53;
   wire multiplier_0_n_54;
   wire multiplier_0_n_55;
   wire multiplier_0_n_56;
   wire multiplier_0_n_57;
   wire multiplier_0_n_136;
   wire multiplier_0_n_119;
   wire multiplier_0_n_69;
   wire multiplier_0_n_121;
   wire multiplier_0_n_88;
   wire multiplier_0_n_90;
   wire multiplier_0_n_135;
   wire multiplier_0_n_118;
   wire multiplier_0_n_91;
   wire multiplier_0_n_134;
   wire multiplier_0_n_117;
   wire multiplier_0_n_92;
   wire multiplier_0_n_133;
   wire multiplier_0_n_116;
   wire multiplier_0_n_93;
   wire multiplier_0_n_44;
   wire multiplier_0_n_132;
   wire multiplier_0_n_115;
   wire multiplier_0_n_94;
   wire multiplier_0_n_43;
   wire multiplier_0_n_131;
   wire multiplier_0_n_114;
   wire multiplier_0_n_95;
   wire multiplier_0_n_42;
   wire multiplier_0_n_130;
   wire multiplier_0_n_113;
   wire multiplier_0_n_96;
   wire multiplier_0_n_129;
   wire multiplier_0_n_112;
   wire multiplier_0_n_97;
   wire multiplier_0_n_128;
   wire multiplier_0_n_111;
   wire multiplier_0_n_98;
   wire multiplier_0_n_127;
   wire multiplier_0_n_110;
   wire multiplier_0_n_99;
   wire multiplier_0_n_126;
   wire multiplier_0_n_109;
   wire multiplier_0_n_100;
   wire multiplier_0_n_125;
   wire multiplier_0_n_108;
   wire multiplier_0_n_101;
   wire multiplier_0_n_124;
   wire multiplier_0_n_107;
   wire multiplier_0_n_102;
   wire multiplier_0_n_123;
   wire multiplier_0_n_106;
   wire multiplier_0_n_103;
   wire multiplier_0_n_122;
   wire multiplier_0_n_105;
   wire multiplier_0_n_104;
   wire multiplier_0_n_89;
   wire multiplier_0_n_137;
   wire multiplier_0_n_120;
   wire multiplier_0_n_0;
   wire multiplier_0_n_13;
   wire multiplier_0_n_9;
   wire multiplier_0_n_11;
   wire multiplier_0_n_10;
   wire multiplier_0_n_150;
   wire multiplier_0_n_58;
   wire multiplier_0_n_59;
   wire multiplier_0_n_60;
   wire multiplier_0_n_61;
   wire multiplier_0_n_62;
   wire multiplier_0_n_63;
   wire multiplier_0_n_64;
   wire multiplier_0_n_65;
   wire multiplier_0_n_66;
   wire multiplier_0_n_7;
   wire multiplier_0_n_86;
   wire multiplier_0_n_87;
   wire multiplier_0_n_70;
   wire multiplier_0_n_85;
   wire multiplier_0_n_84;
   wire multiplier_0_n_83;
   wire multiplier_0_n_82;
   wire multiplier_0_n_81;
   wire multiplier_0_n_80;
   wire multiplier_0_n_79;
   wire multiplier_0_n_78;
   wire multiplier_0_n_77;
   wire multiplier_0_n_76;
   wire multiplier_0_n_75;
   wire multiplier_0_n_74;
   wire multiplier_0_n_73;
   wire multiplier_0_n_72;
   wire multiplier_0_n_71;
   wire multiplier_0_n_138;
   wire multiplier_0_n_142;
   wire multiplier_0_n_143;
   wire multiplier_0_n_140;
   wire multiplier_0_n_148;
   wire multiplier_0_n_8;
   wire multiplier_0_n_149;
   wire multiplier_0_n_12;
   wire multiplier_0_n_37;
   wire multiplier_0_n_14;
   wire multiplier_0_n_36;
   wire multiplier_0_n_35;
   wire multiplier_0_n_34;
   wire multiplier_0_n_33;
   wire multiplier_0_n_32;
   wire multiplier_0_n_31;
   wire multiplier_0_n_30;
   wire multiplier_0_n_29;
   wire multiplier_0_n_28;
   wire multiplier_0_n_27;
   wire multiplier_0_n_26;
   wire multiplier_0_n_25;
   wire multiplier_0_n_24;
   wire multiplier_0_n_145;
   wire multiplier_0_n_147;
   wire multiplier_0_n_23;
   wire multiplier_0_n_139;
   wire multiplier_0_n_141;
   wire multiplier_0_n_144;
   wire multiplier_0_n_146;
   wire multiplier_0_n_22;
   wire mem_backbone_0_n_0_0;
   wire [15:0]mem_backbone_0_per_dout_val;
   wire mem_backbone_0_n_2_0;
   wire mem_backbone_0_n_2_1;
   wire [14:0]mem_backbone_0_ext_mem_addr;
   wire mem_backbone_0_n_2_2;
   wire mem_backbone_0_n_2_3;
   wire mem_backbone_0_n_2_4;
   wire mem_backbone_0_n_2_5;
   wire mem_backbone_0_n_2_6;
   wire mem_backbone_0_n_2_7;
   wire mem_backbone_0_n_2_8;
   wire mem_backbone_0_n_2_9;
   wire mem_backbone_0_n_2_10;
   wire mem_backbone_0_n_2_11;
   wire mem_backbone_0_n_2_12;
   wire mem_backbone_0_n_2_13;
   wire mem_backbone_0_n_2_14;
   wire mem_backbone_0_n_2_15;
   wire mem_backbone_0_n_3_0;
   wire mem_backbone_0_ext_per_sel;
   wire mem_backbone_0_ext_mem_en;
   wire mem_backbone_0_n_5_0;
   wire mem_backbone_0_n_5_1;
   wire mem_backbone_0_n_5_2;
   wire mem_backbone_0_eu_per_en;
   wire mem_backbone_0_n_6_0;
   wire mem_backbone_0_ext_per_en;
   wire mem_backbone_0_ext_pmem_sel;
   wire mem_backbone_0_n_8_0;
   wire mem_backbone_0_fe_pmem_en;
   wire mem_backbone_0_n_11_0;
   wire mem_backbone_0_n_11_1;
   wire mem_backbone_0_eu_pmem_en;
   wire mem_backbone_0_n_12_0;
   wire mem_backbone_0_ext_pmem_en;
   wire [1:0]mem_backbone_0_ext_mem_din_sel;
   wire mem_backbone_0_n_15_0;
   wire mem_backbone_0_n_16_0;
   wire mem_backbone_0_n_16_1;
   wire mem_backbone_0_n_16_2;
   wire mem_backbone_0_n_16_3;
   wire mem_backbone_0_n_16_4;
   wire mem_backbone_0_n_16_5;
   wire mem_backbone_0_n_16_6;
   wire mem_backbone_0_n_16_7;
   wire mem_backbone_0_n_16_8;
   wire mem_backbone_0_n_16_9;
   wire mem_backbone_0_n_16_10;
   wire mem_backbone_0_n_16_11;
   wire mem_backbone_0_n_16_12;
   wire mem_backbone_0_n_16_13;
   wire mem_backbone_0_n_16_14;
   wire mem_backbone_0_n_16_15;
   wire mem_backbone_0_n_19_0;
   wire mem_backbone_0_n_19_1;
   wire mem_backbone_0_n_19_2;
   wire mem_backbone_0_n_19_3;
   wire mem_backbone_0_n_19_4;
   wire mem_backbone_0_n_19_5;
   wire mem_backbone_0_n_19_6;
   wire mem_backbone_0_ext_dmem_sel;
   wire mem_backbone_0_n_20_0;
   wire mem_backbone_0_n_20_1;
   wire mem_backbone_0_n_20_2;
   wire mem_backbone_0_n_20_3;
   wire mem_backbone_0_n_20_4;
   wire mem_backbone_0_n_20_5;
   wire mem_backbone_0_eu_dmem_en;
   wire mem_backbone_0_n_21_0;
   wire mem_backbone_0_ext_dmem_en;
   wire mem_backbone_0_n_22_0;
   wire mem_backbone_0_n_22_1;
   wire mem_backbone_0_n_22_2;
   wire mem_backbone_0_n_22_3;
   wire mem_backbone_0_n_22_4;
   wire mem_backbone_0_n_22_5;
   wire mem_backbone_0_n_22_6;
   wire mem_backbone_0_n_22_7;
   wire mem_backbone_0_n_22_8;
   wire mem_backbone_0_n_22_9;
   wire mem_backbone_0_n_24_0;
   wire mem_backbone_0_n_24_1;
   wire mem_backbone_0_n_24_2;
   wire mem_backbone_0_n_24_3;
   wire mem_backbone_0_n_24_4;
   wire mem_backbone_0_n_24_5;
   wire mem_backbone_0_n_24_6;
   wire mem_backbone_0_n_24_7;
   wire mem_backbone_0_n_24_8;
   wire mem_backbone_0_n_24_9;
   wire mem_backbone_0_n_24_10;
   wire mem_backbone_0_n_24_11;
   wire mem_backbone_0_n_24_12;
   wire mem_backbone_0_n_24_13;
   wire mem_backbone_0_n_24_14;
   wire mem_backbone_0_n_24_15;
   wire mem_backbone_0_n_24_16;
   wire mem_backbone_0_n_25_0;
   wire mem_backbone_0_n_25_1;
   wire mem_backbone_0_n_25_2;
   wire mem_backbone_0_n_25_3;
   wire mem_backbone_0_n_25_4;
   wire mem_backbone_0_n_25_5;
   wire mem_backbone_0_n_25_6;
   wire mem_backbone_0_n_25_7;
   wire mem_backbone_0_n_25_8;
   wire mem_backbone_0_n_25_9;
   wire mem_backbone_0_n_25_10;
   wire mem_backbone_0_n_25_11;
   wire mem_backbone_0_n_25_12;
   wire mem_backbone_0_n_25_13;
   wire mem_backbone_0_n_25_14;
   wire mem_backbone_0_n_25_15;
   wire mem_backbone_0_n_25_16;
   wire mem_backbone_0_n_27_0;
   wire mem_backbone_0_n_27_1;
   wire [1:0]mem_backbone_0_ext_mem_wr;
   wire mem_backbone_0_n_27_2;
   wire mem_backbone_0_n_29_0;
   wire mem_backbone_0_n_29_1;
   wire mem_backbone_0_n_29_2;
   wire [1:0]mem_backbone_0_eu_mdb_in_sel;
   wire mem_backbone_0_n_31_0;
   wire mem_backbone_0_n_32_0;
   wire mem_backbone_0_n_32_1;
   wire mem_backbone_0_n_32_2;
   wire mem_backbone_0_n_32_3;
   wire mem_backbone_0_n_32_4;
   wire mem_backbone_0_n_32_5;
   wire mem_backbone_0_n_32_6;
   wire mem_backbone_0_n_32_7;
   wire mem_backbone_0_n_32_8;
   wire mem_backbone_0_n_32_9;
   wire mem_backbone_0_n_32_10;
   wire mem_backbone_0_n_32_11;
   wire mem_backbone_0_n_32_12;
   wire mem_backbone_0_n_32_13;
   wire mem_backbone_0_n_32_14;
   wire mem_backbone_0_n_32_15;
   wire mem_backbone_0_fe_pmem_en_dly;
   wire mem_backbone_0_n_33_0;
   wire mem_backbone_0_fe_pmem_save;
   wire [15:0]mem_backbone_0_pmem_dout_bckup;
   wire mem_backbone_0_n_35_0;
   wire mem_backbone_0_n_35_1;
   wire mem_backbone_0_fe_pmem_restore;
   wire mem_backbone_0_pmem_dout_bckup_sel;
   wire mem_backbone_0_n_37_0;
   wire mem_backbone_0_n_37_1;
   wire mem_backbone_0_n_39_0;
   wire mem_backbone_0_n_39_1;
   wire mem_backbone_0_n_39_2;
   wire mem_backbone_0_n_39_3;
   wire mem_backbone_0_n_39_4;
   wire mem_backbone_0_n_39_5;
   wire mem_backbone_0_n_39_6;
   wire mem_backbone_0_n_39_7;
   wire mem_backbone_0_n_39_8;
   wire mem_backbone_0_n_39_9;
   wire mem_backbone_0_n_39_10;
   wire mem_backbone_0_n_39_11;
   wire mem_backbone_0_n_39_12;
   wire mem_backbone_0_n_39_13;
   wire mem_backbone_0_n_39_14;
   wire mem_backbone_0_n_39_15;
   wire mem_backbone_0_n_39_16;
   wire mem_backbone_0_n_42_0;
   wire mem_backbone_0_n_43_0;
   wire mem_backbone_0_dma_ready_dly;
   wire mem_backbone_0_n_45_0;
   wire mem_backbone_0_n_45_1;
   wire mem_backbone_0_n_45_2;
   wire mem_backbone_0_n_45_3;
   wire mem_backbone_0_n_45_4;
   wire mem_backbone_0_n_45_5;
   wire mem_backbone_0_n_45_6;
   wire mem_backbone_0_n_45_7;
   wire mem_backbone_0_n_45_8;
   wire mem_backbone_0_n_46_0;
   wire mem_backbone_0_n_46_1;
   wire mem_backbone_0_n_46_2;
   wire mem_backbone_0_n_46_3;
   wire mem_backbone_0_n_46_4;
   wire mem_backbone_0_n_46_5;
   wire mem_backbone_0_n_46_6;
   wire mem_backbone_0_n_46_7;
   wire mem_backbone_0_n_46_8;
   wire mem_backbone_0_n_46_9;
   wire mem_backbone_0_n_46_10;
   wire mem_backbone_0_n_46_11;
   wire mem_backbone_0_n_46_12;
   wire mem_backbone_0_n_46_13;
   wire mem_backbone_0_n_46_14;
   wire mem_backbone_0_n_46_15;
   wire mem_backbone_0_n_46_16;
   wire mem_backbone_0_n_47_0;
   wire mem_backbone_0_n_47_1;
   wire mem_backbone_0_n_47_2;
   wire mem_backbone_0_n_49_0;
   wire mem_backbone_0_n_49_1;
   wire mem_backbone_0_n_49_2;
   wire mem_backbone_0_n_49_3;
   wire mem_backbone_0_n_49_4;
   wire mem_backbone_0_n_49_5;
   wire mem_backbone_0_n_49_6;
   wire mem_backbone_0_n_49_7;
   wire mem_backbone_0_n_49_8;
   wire mem_backbone_0_n_49_9;
   wire mem_backbone_0_n_49_10;
   wire mem_backbone_0_n_49_11;
   wire mem_backbone_0_n_51_0;
   wire mem_backbone_0_n_51_1;
   wire mem_backbone_0_n_0;
   wire mem_backbone_0_n_1;
   wire mem_backbone_0_n_2;
   wire mem_backbone_0_n_4;
   wire mem_backbone_0_n_3;
   wire mem_backbone_0_n_5;
   wire mem_backbone_0_n_6;
   wire mem_backbone_0_n_8;
   wire mem_backbone_0_n_10;
   wire mem_backbone_0_n_7;
   wire mem_backbone_0_n_9;
   wire mem_backbone_0_n_12;
   wire mem_backbone_0_n_11;
   wire mem_backbone_0_n_15;
   wire mem_backbone_0_n_14;
   wire mem_backbone_0_n_13;
   wire mem_backbone_0_n_16;
   wire frontend_0_mirq_wkup;
   wire frontend_0_n_0_0;
   wire frontend_0_cpu_halt_req;
   wire frontend_0_n_3_0;
   wire frontend_0_n_3_1;
   wire frontend_0_n_3_2;
   wire frontend_0_n_3_3;
   wire frontend_0_n_4_0;
   wire frontend_0_n_4_1;
   wire frontend_0_n_4_2;
   wire [2:0]frontend_0_i_state;
   wire frontend_0_n_6_0;
   wire frontend_0_n_6_1;
   wire frontend_0_n_6_2;
   wire frontend_0_n_10_0;
   wire frontend_0_n_10_1;
   wire [3:0]frontend_0_src_reg;
   wire frontend_0_n_10_2;
   wire frontend_0_n_10_3;
   wire frontend_0_n_10_4;
   wire frontend_0_n_11_0;
   wire frontend_0_inst_type_nxt;
   wire frontend_0_n_12_0;
   wire frontend_0_n_12_1;
   wire frontend_0_n_12_2;
   wire frontend_0_n_12_3;
   wire frontend_0_n_12_4;
   wire frontend_0_n_12_5;
   wire frontend_0_n_12_6;
   wire frontend_0_n_12_7;
   wire frontend_0_n_12_8;
   wire frontend_0_n_12_9;
   wire [12:0]frontend_0_inst_as_nxt;
   wire frontend_0_n_12_10;
   wire frontend_0_n_12_11;
   wire frontend_0_n_12_12;
   wire frontend_0_n_12_13;
   wire frontend_0_n_12_14;
   wire frontend_0_n_13_0;
   wire frontend_0_n_13_1;
   wire frontend_0_is_const;
   wire frontend_0_is_sext;
   wire frontend_0_n_16_0;
   wire frontend_0_inst_dext_rdy;
   wire frontend_0_exec_dext_rdy;
   wire frontend_0_n_19_0;
   wire frontend_0_n_19_1;
   wire frontend_0_n_20_0;
   wire frontend_0_n_20_1;
   wire frontend_0_n_20_2;
   wire frontend_0_n_20_3;
   wire frontend_0_n_22_0;
   wire frontend_0_n_23_0;
   wire frontend_0_n_23_1;
   wire frontend_0_n_23_2;
   wire frontend_0_n_23_3;
   wire frontend_0_n_23_4;
   wire frontend_0_n_23_5;
   wire frontend_0_n_23_6;
   wire frontend_0_n_23_7;
   wire frontend_0_n_23_8;
   wire frontend_0_n_23_9;
   wire frontend_0_n_23_10;
   wire frontend_0_n_23_11;
   wire frontend_0_n_23_12;
   wire frontend_0_n_23_13;
   wire frontend_0_n_23_14;
   wire frontend_0_n_23_15;
   wire frontend_0_n_23_16;
   wire frontend_0_n_23_17;
   wire frontend_0_inst_ad_nxt;
   wire frontend_0_n_25_0;
   wire frontend_0_n_25_1;
   wire frontend_0_n_25_2;
   wire frontend_0_n_25_3;
   wire frontend_0_n_25_4;
   wire frontend_0_n_25_5;
   wire frontend_0_n_25_6;
   wire frontend_0_n_27_0;
   wire [7:0]frontend_0_inst_so_nxt;
   wire frontend_0_n_27_1;
   wire frontend_0_inst_sext_rdy;
   wire frontend_0_exec_dst_wr;
   wire frontend_0_n_32_0;
   wire frontend_0_n_33_0;
   wire frontend_0_n_33_1;
   wire frontend_0_n_33_2;
   wire frontend_0_n_33_3;
   wire frontend_0_n_33_4;
   wire frontend_0_exec_src_wr;
   wire frontend_0_n_39_0;
   wire frontend_0_n_39_1;
   wire frontend_0_exec_jmp;
   wire frontend_0_n_44_0;
   wire frontend_0_n_44_1;
   wire frontend_0_n_45_0;
   wire frontend_0_n_45_1;
   wire frontend_0_n_45_2;
   wire frontend_0_dst_acalc_pre;
   wire frontend_0_src_acalc_pre;
   wire frontend_0_n_50_0;
   wire frontend_0_n_50_1;
   wire frontend_0_n_50_2;
   wire frontend_0_n_50_3;
   wire frontend_0_n_50_4;
   wire frontend_0_n_50_5;
   wire frontend_0_n_50_6;
   wire frontend_0_n_50_7;
   wire frontend_0_n_50_8;
   wire frontend_0_n_50_9;
   wire frontend_0_n_50_10;
   wire frontend_0_n_50_11;
   wire frontend_0_n_50_12;
   wire frontend_0_n_50_13;
   wire frontend_0_n_50_14;
   wire frontend_0_n_50_15;
   wire frontend_0_n_50_16;
   wire frontend_0_n_50_17;
   wire frontend_0_n_50_18;
   wire frontend_0_n_50_19;
   wire frontend_0_n_53_0;
   wire frontend_0_n_53_1;
   wire frontend_0_n_55_0;
   wire frontend_0_n_55_1;
   wire frontend_0_n_55_2;
   wire frontend_0_n_55_3;
   wire frontend_0_n_55_4;
   wire frontend_0_n_55_5;
   wire frontend_0_n_55_6;
   wire frontend_0_n_55_7;
   wire frontend_0_n_55_8;
   wire frontend_0_n_55_9;
   wire frontend_0_n_55_10;
   wire frontend_0_n_55_11;
   wire frontend_0_n_55_12;
   wire frontend_0_n_55_13;
   wire frontend_0_n_55_14;
   wire frontend_0_n_55_15;
   wire frontend_0_n_55_16;
   wire frontend_0_n_55_17;
   wire frontend_0_n_55_18;
   wire frontend_0_n_55_19;
   wire frontend_0_n_55_20;
   wire frontend_0_n_55_21;
   wire frontend_0_n_55_22;
   wire frontend_0_n_55_23;
   wire frontend_0_n_55_24;
   wire frontend_0_n_55_25;
   wire frontend_0_n_55_26;
   wire frontend_0_n_55_27;
   wire frontend_0_n_55_28;
   wire frontend_0_n_55_29;
   wire frontend_0_n_55_30;
   wire frontend_0_n_55_31;
   wire frontend_0_n_55_32;
   wire frontend_0_n_55_33;
   wire frontend_0_n_55_34;
   wire [3:0]frontend_0_e_state_nxt_reg;
   wire frontend_0_n_55_35;
   wire frontend_0_n_55_36;
   wire frontend_0_n_55_37;
   wire frontend_0_n_55_38;
   wire frontend_0_n_55_39;
   wire frontend_0_n_55_40;
   wire frontend_0_n_55_41;
   wire frontend_0_n_55_42;
   wire frontend_0_n_55_43;
   wire frontend_0_n_55_44;
   wire frontend_0_n_55_45;
   wire frontend_0_n_55_46;
   wire frontend_0_n_55_47;
   wire frontend_0_n_55_48;
   wire frontend_0_n_55_49;
   wire frontend_0_n_55_50;
   wire frontend_0_n_55_51;
   wire frontend_0_n_55_52;
   wire frontend_0_n_55_53;
   wire frontend_0_n_55_54;
   wire frontend_0_n_55_55;
   wire frontend_0_n_55_56;
   wire frontend_0_n_55_57;
   wire frontend_0_n_55_58;
   wire frontend_0_n_55_59;
   wire frontend_0_n_55_60;
   wire frontend_0_n_55_61;
   wire frontend_0_n_55_62;
   wire frontend_0_n_55_63;
   wire frontend_0_n_55_64;
   wire frontend_0_n_55_65;
   wire frontend_0_n_55_66;
   wire frontend_0_n_55_67;
   wire frontend_0_n_55_68;
   wire frontend_0_n_58_0;
   wire frontend_0_n_58_1;
   wire frontend_0_n_58_2;
   wire frontend_0_n_58_3;
   wire frontend_0_n_59_0;
   wire frontend_0_n_59_1;
   wire frontend_0_n_59_2;
   wire frontend_0_n_59_3;
   wire frontend_0_n_59_4;
   wire frontend_0_n_59_5;
   wire frontend_0_n_59_6;
   wire frontend_0_n_60_0;
   wire frontend_0_irq_detect;
   wire frontend_0_decode;
   wire frontend_0_n_64_0;
   wire [1:0]frontend_0_inst_sz_nxt;
   wire [1:0]frontend_0_inst_sz;
   wire frontend_0_n_70_0;
   wire frontend_0_n_71_0;
   wire frontend_0_n_72_0;
   wire frontend_0_n_73_0;
   wire frontend_0_n_73_1;
   wire frontend_0_n_73_2;
   wire frontend_0_n_73_3;
   wire frontend_0_n_74_0;
   wire frontend_0_n_75_0;
   wire frontend_0_n_76_0;
   wire frontend_0_n_76_1;
   wire frontend_0_n_76_2;
   wire frontend_0_n_76_3;
   wire frontend_0_n_76_4;
   wire frontend_0_n_76_5;
   wire frontend_0_n_76_6;
   wire frontend_0_n_76_7;
   wire [2:0]frontend_0_i_state_nxt_reg;
   wire frontend_0_n_76_8;
   wire frontend_0_n_76_9;
   wire frontend_0_n_76_10;
   wire frontend_0_n_76_11;
   wire frontend_0_n_76_12;
   wire frontend_0_n_76_13;
   wire frontend_0_n_76_14;
   wire frontend_0_n_80_0;
   wire frontend_0_n_82_0;
   wire frontend_0_n_82_1;
   wire frontend_0_n_82_2;
   wire frontend_0_n_82_3;
   wire frontend_0_n_82_4;
   wire frontend_0_n_82_5;
   wire frontend_0_n_82_6;
   wire frontend_0_n_82_7;
   wire frontend_0_n_82_8;
   wire frontend_0_n_82_9;
   wire frontend_0_n_82_10;
   wire [11:0]frontend_0_inst_to_nxt;
   wire frontend_0_alu_inc;
   wire [11:0]frontend_0_inst_alu_nxt;
   wire frontend_0_n_88_0;
   wire frontend_0_n_88_1;
   wire frontend_0_n_91_0;
   wire [3:0]frontend_0_inst_dest_bin;
   wire frontend_0_n_94_0;
   wire frontend_0_n_94_1;
   wire frontend_0_n_94_2;
   wire frontend_0_n_94_3;
   wire frontend_0_n_94_4;
   wire frontend_0_n_94_5;
   wire frontend_0_n_94_6;
   wire frontend_0_n_94_7;
   wire frontend_0_n_94_8;
   wire frontend_0_n_94_9;
   wire frontend_0_n_94_10;
   wire frontend_0_n_94_11;
   wire frontend_0_n_95_0;
   wire frontend_0_n_95_1;
   wire frontend_0_n_95_2;
   wire frontend_0_n_95_3;
   wire frontend_0_n_95_4;
   wire frontend_0_n_95_5;
   wire frontend_0_n_95_6;
   wire frontend_0_n_95_7;
   wire frontend_0_n_95_8;
   wire frontend_0_n_95_9;
   wire frontend_0_n_95_10;
   wire frontend_0_n_95_11;
   wire frontend_0_n_97_0;
   wire frontend_0_n_97_1;
   wire frontend_0_n_97_2;
   wire frontend_0_n_97_3;
   wire frontend_0_n_97_4;
   wire frontend_0_n_97_5;
   wire frontend_0_n_97_6;
   wire frontend_0_n_97_7;
   wire frontend_0_n_97_8;
   wire frontend_0_n_97_9;
   wire frontend_0_n_97_10;
   wire frontend_0_n_97_11;
   wire frontend_0_n_97_12;
   wire frontend_0_n_97_13;
   wire frontend_0_n_97_14;
   wire frontend_0_n_97_15;
   wire frontend_0_n_97_16;
   wire frontend_0_n_97_17;
   wire frontend_0_n_97_18;
   wire frontend_0_n_97_19;
   wire frontend_0_n_98_0;
   wire frontend_0_n_98_1;
   wire frontend_0_n_98_2;
   wire frontend_0_n_98_3;
   wire frontend_0_n_98_4;
   wire frontend_0_n_99_0;
   wire [15:0]frontend_0_ext_nxt;
   wire frontend_0_n_99_1;
   wire frontend_0_n_99_2;
   wire frontend_0_n_99_3;
   wire frontend_0_n_99_4;
   wire frontend_0_n_99_5;
   wire frontend_0_n_99_6;
   wire frontend_0_n_99_7;
   wire frontend_0_n_99_8;
   wire frontend_0_n_99_9;
   wire frontend_0_n_99_10;
   wire frontend_0_n_99_11;
   wire frontend_0_n_99_12;
   wire frontend_0_n_99_13;
   wire frontend_0_n_99_14;
   wire frontend_0_n_99_15;
   wire frontend_0_n_99_16;
   wire frontend_0_n_99_17;
   wire frontend_0_n_101_0;
   wire frontend_0_n_101_1;
   wire [2:0]frontend_0_inst_jmp_bin;
   wire frontend_0_n_105_0;
   wire frontend_0_n_105_1;
   wire frontend_0_n_105_2;
   wire frontend_0_n_105_3;
   wire frontend_0_n_105_4;
   wire frontend_0_n_105_5;
   wire frontend_0_n_105_6;
   wire frontend_0_n_110_0;
   wire frontend_0_n_110_1;
   wire frontend_0_n_110_2;
   wire frontend_0_n_110_3;
   wire frontend_0_n_110_4;
   wire frontend_0_n_110_5;
   wire frontend_0_n_110_6;
   wire frontend_0_n_110_7;
   wire frontend_0_n_110_8;
   wire frontend_0_n_110_9;
   wire frontend_0_n_110_10;
   wire frontend_0_n_110_11;
   wire frontend_0_n_110_12;
   wire frontend_0_n_110_13;
   wire frontend_0_n_110_14;
   wire frontend_0_n_110_15;
   wire frontend_0_n_110_16;
   wire frontend_0_n_110_17;
   wire frontend_0_n_110_18;
   wire frontend_0_n_110_19;
   wire frontend_0_n_110_20;
   wire frontend_0_n_110_21;
   wire frontend_0_n_110_22;
   wire frontend_0_n_110_23;
   wire frontend_0_n_110_24;
   wire frontend_0_n_110_25;
   wire frontend_0_n_110_26;
   wire frontend_0_n_110_27;
   wire frontend_0_n_110_28;
   wire frontend_0_n_110_29;
   wire frontend_0_n_110_30;
   wire frontend_0_n_110_31;
   wire frontend_0_n_110_32;
   wire frontend_0_n_110_33;
   wire frontend_0_n_110_34;
   wire frontend_0_n_110_35;
   wire frontend_0_n_111_0;
   wire frontend_0_n_111_1;
   wire frontend_0_n_111_2;
   wire frontend_0_n_111_3;
   wire frontend_0_n_111_4;
   wire [3:0]frontend_0_inst_src_bin;
   wire frontend_0_n_114_0;
   wire frontend_0_n_114_1;
   wire frontend_0_n_114_2;
   wire frontend_0_n_114_3;
   wire frontend_0_n_114_4;
   wire frontend_0_n_114_5;
   wire frontend_0_n_114_6;
   wire frontend_0_n_114_7;
   wire frontend_0_n_114_8;
   wire frontend_0_n_114_9;
   wire frontend_0_n_114_10;
   wire frontend_0_n_114_11;
   wire frontend_0_n_115_0;
   wire frontend_0_n_115_1;
   wire frontend_0_n_115_2;
   wire frontend_0_n_115_3;
   wire frontend_0_n_115_4;
   wire frontend_0_n_115_5;
   wire frontend_0_n_115_6;
   wire frontend_0_n_115_7;
   wire frontend_0_n_115_8;
   wire frontend_0_n_115_9;
   wire frontend_0_n_115_10;
   wire frontend_0_n_115_11;
   wire frontend_0_n_115_12;
   wire frontend_0_n_115_13;
   wire frontend_0_n_115_14;
   wire frontend_0_n_115_15;
   wire frontend_0_n_115_16;
   wire frontend_0_n_115_17;
   wire frontend_0_n_115_18;
   wire frontend_0_n_115_19;
   wire [5:0]frontend_0_irq_num;
   wire frontend_0_n_118_0;
   wire frontend_0_n_118_1;
   wire frontend_0_n_118_2;
   wire frontend_0_n_118_3;
   wire frontend_0_n_118_4;
   wire frontend_0_n_118_5;
   wire frontend_0_n_118_6;
   wire frontend_0_n_118_7;
   wire frontend_0_n_118_8;
   wire frontend_0_n_118_9;
   wire frontend_0_n_118_10;
   wire frontend_0_n_118_11;
   wire frontend_0_n_118_12;
   wire frontend_0_n_118_13;
   wire frontend_0_n_118_14;
   wire frontend_0_n_118_15;
   wire frontend_0_n_118_16;
   wire frontend_0_n_118_17;
   wire frontend_0_n_118_18;
   wire frontend_0_n_118_19;
   wire frontend_0_n_118_20;
   wire frontend_0_n_118_21;
   wire frontend_0_n_118_22;
   wire frontend_0_n_118_23;
   wire frontend_0_n_118_24;
   wire frontend_0_n_118_25;
   wire frontend_0_n_118_26;
   wire frontend_0_n_118_27;
   wire frontend_0_n_118_28;
   wire frontend_0_n_118_29;
   wire frontend_0_n_118_30;
   wire frontend_0_n_118_31;
   wire frontend_0_n_118_32;
   wire frontend_0_n_118_33;
   wire frontend_0_n_118_34;
   wire frontend_0_n_118_35;
   wire frontend_0_n_118_36;
   wire frontend_0_n_118_37;
   wire frontend_0_n_118_38;
   wire frontend_0_n_118_39;
   wire frontend_0_n_118_40;
   wire frontend_0_n_118_41;
   wire frontend_0_n_118_42;
   wire frontend_0_n_118_43;
   wire frontend_0_n_118_44;
   wire frontend_0_n_118_45;
   wire frontend_0_n_118_46;
   wire frontend_0_n_118_47;
   wire frontend_0_n_118_48;
   wire frontend_0_n_118_49;
   wire frontend_0_n_118_50;
   wire frontend_0_n_118_51;
   wire frontend_0_n_118_52;
   wire frontend_0_n_118_53;
   wire frontend_0_n_118_54;
   wire frontend_0_n_118_55;
   wire frontend_0_n_118_56;
   wire frontend_0_n_120_0;
   wire frontend_0_n_120_1;
   wire frontend_0_n_120_2;
   wire frontend_0_n_120_3;
   wire frontend_0_n_120_4;
   wire frontend_0_n_120_5;
   wire frontend_0_n_120_6;
   wire frontend_0_n_120_7;
   wire frontend_0_n_120_8;
   wire frontend_0_n_120_9;
   wire frontend_0_n_120_10;
   wire frontend_0_n_120_11;
   wire frontend_0_n_120_12;
   wire frontend_0_n_120_13;
   wire frontend_0_n_120_14;
   wire frontend_0_n_120_15;
   wire frontend_0_n_120_16;
   wire frontend_0_n_120_17;
   wire frontend_0_n_120_18;
   wire frontend_0_n_120_19;
   wire frontend_0_n_120_20;
   wire frontend_0_n_122_0;
   wire frontend_0_n_122_1;
   wire frontend_0_n_122_2;
   wire frontend_0_fetch;
   wire [15:0]frontend_0_pc_incr;
   wire frontend_0_n_124_0;
   wire frontend_0_n_124_1;
   wire frontend_0_n_124_2;
   wire frontend_0_n_124_3;
   wire frontend_0_n_124_4;
   wire frontend_0_n_124_5;
   wire frontend_0_n_124_6;
   wire frontend_0_n_124_7;
   wire frontend_0_n_124_8;
   wire frontend_0_n_124_9;
   wire frontend_0_n_124_10;
   wire frontend_0_n_124_11;
   wire frontend_0_n_124_12;
   wire frontend_0_n_124_13;
   wire frontend_0_n_124_14;
   wire frontend_0_n_125_0;
   wire frontend_0_n_126_0;
   wire frontend_0_n_126_1;
   wire frontend_0_n_126_2;
   wire frontend_0_n_126_3;
   wire frontend_0_n_126_4;
   wire frontend_0_n_126_5;
   wire frontend_0_n_126_6;
   wire frontend_0_n_126_7;
   wire frontend_0_n_126_8;
   wire frontend_0_n_126_9;
   wire frontend_0_n_126_10;
   wire frontend_0_n_126_11;
   wire frontend_0_n_126_12;
   wire frontend_0_n_126_13;
   wire frontend_0_n_126_14;
   wire frontend_0_n_126_15;
   wire frontend_0_n_127_0;
   wire frontend_0_n_127_1;
   wire frontend_0_n_127_2;
   wire frontend_0_n_127_3;
   wire frontend_0_n_127_4;
   wire frontend_0_n_127_5;
   wire frontend_0_n_127_6;
   wire frontend_0_n_127_7;
   wire frontend_0_n_127_8;
   wire frontend_0_n_127_9;
   wire frontend_0_n_127_10;
   wire frontend_0_n_127_11;
   wire frontend_0_n_127_12;
   wire frontend_0_n_127_13;
   wire frontend_0_n_127_14;
   wire frontend_0_n_127_15;
   wire frontend_0_n_127_16;
   wire frontend_0_pmem_busy;
   wire frontend_0_n_128_0;
   wire frontend_0_n_128_1;
   wire frontend_0_n_130_0;
   wire frontend_0_n_130_1;
   wire frontend_0_n_130_2;
   wire frontend_0_n_130_3;
   wire frontend_0_n_91;
   wire frontend_0_n_0;
   wire frontend_0_n_87;
   wire frontend_0_n_1;
   wire frontend_0_n_2;
   wire frontend_0_n_3;
   wire frontend_0_n_88;
   wire frontend_0_n_89;
   wire frontend_0_n_5;
   wire frontend_0_n_55;
   wire frontend_0_n_10;
   wire frontend_0_n_29;
   wire frontend_0_n_37;
   wire frontend_0_n_28;
   wire frontend_0_n_36;
   wire frontend_0_n_9;
   wire frontend_0_n_49;
   wire frontend_0_n_17;
   wire frontend_0_n_18;
   wire frontend_0_n_48;
   wire frontend_0_n_4;
   wire frontend_0_n_67;
   wire frontend_0_n_73;
   wire frontend_0_n_51;
   wire frontend_0_n_52;
   wire frontend_0_n_50;
   wire frontend_0_n_11;
   wire frontend_0_n_43;
   wire frontend_0_n_68;
   wire frontend_0_n_45;
   wire frontend_0_n_69;
   wire frontend_0_n_70;
   wire frontend_0_n_46;
   wire frontend_0_n_47;
   wire frontend_0_n_44;
   wire frontend_0_n_72;
   wire frontend_0_n_71;
   wire frontend_0_n_56;
   wire frontend_0_n_54;
   wire frontend_0_n_20;
   wire frontend_0_n_19;
   wire frontend_0_n_26;
   wire frontend_0_n_34;
   wire frontend_0_n_27;
   wire frontend_0_n_35;
   wire frontend_0_n_53;
   wire frontend_0_n_58;
   wire frontend_0_n_6;
   wire frontend_0_n_12;
   wire frontend_0_n_38;
   wire frontend_0_n_39;
   wire frontend_0_n_62;
   wire frontend_0_n_21;
   wire frontend_0_n_63;
   wire frontend_0_n_64;
   wire frontend_0_n_57;
   wire frontend_0_n_13;
   wire frontend_0_n_7;
   wire frontend_0_n_15;
   wire frontend_0_n_16;
   wire frontend_0_n_14;
   wire frontend_0_n_61;
   wire frontend_0_n_66;
   wire frontend_0_n_65;
   wire frontend_0_n_41;
   wire frontend_0_n_42;
   wire frontend_0_n_40;
   wire frontend_0_n_59;
   wire frontend_0_n_60;
   wire frontend_0_n_82;
   wire frontend_0_n_83;
   wire frontend_0_n_86;
   wire frontend_0_n_74;
   wire frontend_0_n_75;
   wire frontend_0_n_76;
   wire frontend_0_n_79;
   wire frontend_0_n_80;
   wire frontend_0_n_90;
   wire frontend_0_n_85;
   wire frontend_0_n_81;
   wire frontend_0_n_77;
   wire frontend_0_n_78;
   wire frontend_0_n_84;
   wire frontend_0_n_92;
   wire frontend_0_n_98;
   wire frontend_0_n_100;
   wire frontend_0_n_108;
   wire frontend_0_n_24;
   wire frontend_0_n_32;
   wire frontend_0_n_22;
   wire frontend_0_n_30;
   wire frontend_0_n_104;
   wire frontend_0_n_107;
   wire frontend_0_n_25;
   wire frontend_0_n_33;
   wire frontend_0_n_94;
   wire frontend_0_n_97;
   wire frontend_0_n_96;
   wire frontend_0_n_95;
   wire frontend_0_n_105;
   wire frontend_0_n_106;
   wire frontend_0_n_103;
   wire frontend_0_n_99;
   wire frontend_0_n_102;
   wire frontend_0_n_101;
   wire frontend_0_n_110;
   wire frontend_0_n_109;
   wire frontend_0_n_144;
   wire frontend_0_n_111;
   wire frontend_0_n_127;
   wire frontend_0_n_143;
   wire frontend_0_n_126;
   wire frontend_0_n_142;
   wire frontend_0_n_125;
   wire frontend_0_n_141;
   wire frontend_0_n_124;
   wire frontend_0_n_140;
   wire frontend_0_n_123;
   wire frontend_0_n_139;
   wire frontend_0_n_122;
   wire frontend_0_n_138;
   wire frontend_0_n_121;
   wire frontend_0_n_137;
   wire frontend_0_n_120;
   wire frontend_0_n_136;
   wire frontend_0_n_119;
   wire frontend_0_n_135;
   wire frontend_0_n_118;
   wire frontend_0_n_134;
   wire frontend_0_n_117;
   wire frontend_0_n_133;
   wire frontend_0_n_116;
   wire frontend_0_n_132;
   wire frontend_0_n_115;
   wire frontend_0_n_131;
   wire frontend_0_n_114;
   wire frontend_0_n_130;
   wire frontend_0_n_113;
   wire frontend_0_n_129;
   wire frontend_0_n_112;
   wire frontend_0_n_128;
   wire frontend_0_n_145;
   wire frontend_0_n_147;
   wire frontend_0_n_146;
   wire frontend_0_n_148;
   wire frontend_0_n_149;
   wire frontend_0_n_157;
   wire frontend_0_n_156;
   wire frontend_0_n_155;
   wire frontend_0_n_154;
   wire frontend_0_n_153;
   wire frontend_0_n_152;
   wire frontend_0_n_151;
   wire frontend_0_n_150;
   wire frontend_0_n_93;
   wire frontend_0_n_158;
   wire frontend_0_n_179;
   wire frontend_0_n_180;
   wire frontend_0_n_163;
   wire frontend_0_n_178;
   wire frontend_0_n_177;
   wire frontend_0_n_176;
   wire frontend_0_n_175;
   wire frontend_0_n_174;
   wire frontend_0_n_173;
   wire frontend_0_n_172;
   wire frontend_0_n_171;
   wire frontend_0_n_170;
   wire frontend_0_n_169;
   wire frontend_0_n_168;
   wire frontend_0_n_162;
   wire frontend_0_n_167;
   wire frontend_0_n_161;
   wire frontend_0_n_166;
   wire frontend_0_n_160;
   wire frontend_0_n_165;
   wire frontend_0_n_159;
   wire frontend_0_n_164;
   wire frontend_0_n_23;
   wire frontend_0_n_31;
   wire frontend_0_n_181;
   wire frontend_0_n_197;
   wire frontend_0_n_196;
   wire frontend_0_n_195;
   wire frontend_0_n_194;
   wire frontend_0_n_193;
   wire frontend_0_n_192;
   wire frontend_0_n_191;
   wire frontend_0_n_190;
   wire frontend_0_n_189;
   wire frontend_0_n_188;
   wire frontend_0_n_187;
   wire frontend_0_n_186;
   wire frontend_0_n_185;
   wire frontend_0_n_184;
   wire frontend_0_n_183;
   wire frontend_0_n_182;
   wire frontend_0_n_8;
   wire frontend_0_n_198;
   wire frontend_0_n_200;
   wire frontend_0_n_199;
   wire frontend_0_n_201;
   wire frontend_0_n_202;
   wire frontend_0_n_203;
   wire frontend_0_n_204;
   wire frontend_0_n_218;
   wire frontend_0_n_217;
   wire frontend_0_n_216;
   wire frontend_0_n_215;
   wire frontend_0_n_214;
   wire frontend_0_n_213;
   wire frontend_0_n_212;
   wire frontend_0_n_211;
   wire frontend_0_n_210;
   wire frontend_0_n_209;
   wire frontend_0_n_208;
   wire frontend_0_n_207;
   wire frontend_0_n_206;
   wire frontend_0_n_205;
   wire frontend_0_n_221;
   wire frontend_0_n_220;
   wire frontend_0_n_222;
   wire frontend_0_n_237;
   wire frontend_0_n_236;
   wire frontend_0_n_235;
   wire frontend_0_n_234;
   wire frontend_0_n_233;
   wire frontend_0_n_232;
   wire frontend_0_n_231;
   wire frontend_0_n_230;
   wire frontend_0_n_229;
   wire frontend_0_n_228;
   wire frontend_0_n_227;
   wire frontend_0_n_226;
   wire frontend_0_n_225;
   wire frontend_0_n_224;
   wire frontend_0_n_238;
   wire frontend_0_n_223;
   wire frontend_0_n_240;
   wire frontend_0_n_239;
   wire frontend_0_n_219;
   wire [3:0]execution_unit_0_alu_stat_wr;
   wire [3:0]execution_unit_0_alu_stat;
   wire [15:0]execution_unit_0_alu_out;
   wire [3:0]execution_unit_0_status;
   wire [15:0]execution_unit_0_reg_src;
   wire execution_unit_0_n_0_0;
   wire execution_unit_0_n_0_1;
   wire execution_unit_0_n_0_2;
   wire execution_unit_0_n_0_3;
   wire execution_unit_0_reg_sr_clr;
   wire execution_unit_0_n_4_0;
   wire execution_unit_0_n_4_1;
   wire execution_unit_0_mb_wr_det;
   wire execution_unit_0_n_7_0;
   wire execution_unit_0_n_7_1;
   wire execution_unit_0_n_7_2;
   wire execution_unit_0_n_7_3;
   wire execution_unit_0_n_7_4;
   wire execution_unit_0_n_8_0;
   wire execution_unit_0_n_8_1;
   wire execution_unit_0_n_8_2;
   wire execution_unit_0_n_8_3;
   wire execution_unit_0_mab_lsb;
   wire [15:0]execution_unit_0_mdb_out_nxt;
   wire execution_unit_0_n_13_0;
   wire execution_unit_0_n_13_1;
   wire execution_unit_0_n_13_2;
   wire execution_unit_0_n_13_3;
   wire execution_unit_0_n_13_4;
   wire execution_unit_0_n_13_5;
   wire execution_unit_0_n_13_6;
   wire execution_unit_0_n_13_7;
   wire execution_unit_0_n_13_8;
   wire execution_unit_0_n_13_9;
   wire execution_unit_0_n_13_10;
   wire execution_unit_0_n_13_11;
   wire execution_unit_0_n_13_12;
   wire execution_unit_0_n_13_13;
   wire execution_unit_0_n_13_14;
   wire execution_unit_0_n_13_15;
   wire execution_unit_0_n_13_16;
   wire execution_unit_0_n_13_17;
   wire execution_unit_0_n_13_18;
   wire execution_unit_0_n_14_0;
   wire execution_unit_0_n_14_1;
   wire execution_unit_0_n_15_0;
   wire execution_unit_0_n_15_1;
   wire execution_unit_0_n_15_2;
   wire execution_unit_0_n_15_3;
   wire execution_unit_0_n_17_0;
   wire execution_unit_0_n_17_1;
   wire execution_unit_0_n_17_2;
   wire execution_unit_0_n_17_3;
   wire execution_unit_0_n_17_4;
   wire execution_unit_0_n_17_5;
   wire execution_unit_0_n_17_6;
   wire execution_unit_0_n_17_7;
   wire execution_unit_0_n_17_8;
   wire execution_unit_0_n_21_0;
   wire execution_unit_0_n_21_1;
   wire execution_unit_0_n_21_2;
   wire execution_unit_0_n_21_3;
   wire execution_unit_0_n_21_4;
   wire execution_unit_0_reg_dest_wr;
   wire execution_unit_0_n_23_0;
   wire execution_unit_0_reg_pc_call;
   wire execution_unit_0_n_30_0;
   wire execution_unit_0_n_30_1;
   wire execution_unit_0_n_30_2;
   wire execution_unit_0_reg_sp_wr;
   wire execution_unit_0_reg_sr_wr;
   wire execution_unit_0_n_32_0;
   wire execution_unit_0_reg_incr;
   wire execution_unit_0_n_34_0;
   wire execution_unit_0_n_34_1;
   wire execution_unit_0_n_34_2;
   wire execution_unit_0_n_34_3;
   wire execution_unit_0_n_34_4;
   wire execution_unit_0_n_34_5;
   wire execution_unit_0_n_34_6;
   wire execution_unit_0_n_34_7;
   wire execution_unit_0_n_34_8;
   wire execution_unit_0_n_34_9;
   wire execution_unit_0_n_34_10;
   wire execution_unit_0_n_34_11;
   wire execution_unit_0_n_34_12;
   wire execution_unit_0_n_34_13;
   wire execution_unit_0_n_34_14;
   wire execution_unit_0_n_34_15;
   wire execution_unit_0_n_34_16;
   wire execution_unit_0_n_34_17;
   wire execution_unit_0_n_39_0;
   wire execution_unit_0_n_39_1;
   wire execution_unit_0_n_39_2;
   wire execution_unit_0_n_39_3;
   wire execution_unit_0_n_39_4;
   wire execution_unit_0_n_39_5;
   wire execution_unit_0_n_39_6;
   wire execution_unit_0_n_39_7;
   wire execution_unit_0_n_39_8;
   wire execution_unit_0_n_40_0;
   wire execution_unit_0_n_40_1;
   wire execution_unit_0_n_40_2;
   wire execution_unit_0_n_40_3;
   wire execution_unit_0_n_40_4;
   wire execution_unit_0_n_40_5;
   wire execution_unit_0_n_40_6;
   wire execution_unit_0_n_41_0;
   wire execution_unit_0_n_41_1;
   wire execution_unit_0_n_41_2;
   wire execution_unit_0_n_41_3;
   wire execution_unit_0_n_41_4;
   wire execution_unit_0_n_41_5;
   wire execution_unit_0_n_41_6;
   wire execution_unit_0_n_41_7;
   wire execution_unit_0_n_41_8;
   wire execution_unit_0_n_41_9;
   wire execution_unit_0_n_41_10;
   wire execution_unit_0_n_41_11;
   wire execution_unit_0_n_41_12;
   wire execution_unit_0_n_41_13;
   wire execution_unit_0_n_41_14;
   wire execution_unit_0_n_41_15;
   wire execution_unit_0_n_41_16;
   wire execution_unit_0_n_41_17;
   wire execution_unit_0_n_41_18;
   wire execution_unit_0_n_41_19;
   wire execution_unit_0_n_41_20;
   wire execution_unit_0_n_41_21;
   wire execution_unit_0_n_41_22;
   wire execution_unit_0_n_41_23;
   wire execution_unit_0_n_41_24;
   wire execution_unit_0_n_41_25;
   wire execution_unit_0_n_41_26;
   wire execution_unit_0_n_41_27;
   wire execution_unit_0_n_41_28;
   wire execution_unit_0_n_41_29;
   wire execution_unit_0_n_41_30;
   wire execution_unit_0_n_41_31;
   wire execution_unit_0_n_41_32;
   wire execution_unit_0_n_41_33;
   wire execution_unit_0_n_41_34;
   wire execution_unit_0_n_41_35;
   wire execution_unit_0_n_41_36;
   wire execution_unit_0_n_41_37;
   wire execution_unit_0_n_41_38;
   wire execution_unit_0_n_41_39;
   wire execution_unit_0_n_41_40;
   wire execution_unit_0_n_41_41;
   wire execution_unit_0_n_41_42;
   wire execution_unit_0_n_41_43;
   wire execution_unit_0_n_41_44;
   wire execution_unit_0_n_41_45;
   wire execution_unit_0_n_41_46;
   wire execution_unit_0_n_41_47;
   wire execution_unit_0_n_41_48;
   wire execution_unit_0_n_41_49;
   wire execution_unit_0_n_41_50;
   wire execution_unit_0_n_41_51;
   wire execution_unit_0_n_41_52;
   wire execution_unit_0_n_41_53;
   wire execution_unit_0_n_41_54;
   wire execution_unit_0_n_41_55;
   wire execution_unit_0_n_41_56;
   wire execution_unit_0_n_41_57;
   wire execution_unit_0_n_41_58;
   wire execution_unit_0_n_41_59;
   wire execution_unit_0_n_41_60;
   wire execution_unit_0_n_41_61;
   wire execution_unit_0_n_41_62;
   wire execution_unit_0_n_41_63;
   wire execution_unit_0_n_41_64;
   wire execution_unit_0_n_41_65;
   wire execution_unit_0_n_41_66;
   wire execution_unit_0_n_41_67;
   wire execution_unit_0_n_41_68;
   wire execution_unit_0_n_41_69;
   wire execution_unit_0_n_41_70;
   wire execution_unit_0_n_41_71;
   wire execution_unit_0_n_41_72;
   wire execution_unit_0_n_41_73;
   wire execution_unit_0_n_41_74;
   wire execution_unit_0_n_41_75;
   wire execution_unit_0_n_41_76;
   wire execution_unit_0_n_41_77;
   wire execution_unit_0_n_41_78;
   wire execution_unit_0_n_41_79;
   wire execution_unit_0_mdb_in_buf_en;
   wire [15:0]execution_unit_0_mdb_in_buf;
   wire execution_unit_0_mdb_in_buf_valid;
   wire execution_unit_0_n_44_0;
   wire execution_unit_0_n_44_1;
   wire execution_unit_0_n_45_0;
   wire execution_unit_0_n_45_1;
   wire execution_unit_0_n_45_2;
   wire execution_unit_0_n_48_0;
   wire execution_unit_0_n_48_1;
   wire execution_unit_0_n_48_2;
   wire execution_unit_0_n_48_3;
   wire execution_unit_0_n_48_4;
   wire execution_unit_0_n_48_5;
   wire execution_unit_0_n_48_6;
   wire execution_unit_0_n_48_7;
   wire execution_unit_0_n_48_8;
   wire execution_unit_0_n_48_9;
   wire execution_unit_0_n_49_0;
   wire execution_unit_0_n_49_1;
   wire execution_unit_0_n_49_2;
   wire execution_unit_0_n_49_3;
   wire execution_unit_0_n_49_4;
   wire execution_unit_0_n_49_5;
   wire execution_unit_0_n_49_6;
   wire execution_unit_0_n_49_7;
   wire execution_unit_0_n_49_8;
   wire execution_unit_0_n_49_9;
   wire execution_unit_0_n_50_0;
   wire execution_unit_0_n_50_1;
   wire execution_unit_0_n_50_2;
   wire execution_unit_0_n_50_3;
   wire execution_unit_0_n_50_4;
   wire execution_unit_0_n_50_5;
   wire execution_unit_0_n_50_6;
   wire execution_unit_0_n_50_7;
   wire execution_unit_0_n_50_8;
   wire execution_unit_0_n_50_9;
   wire execution_unit_0_n_50_10;
   wire execution_unit_0_n_50_11;
   wire execution_unit_0_n_50_12;
   wire execution_unit_0_n_50_13;
   wire execution_unit_0_n_50_14;
   wire execution_unit_0_n_50_15;
   wire execution_unit_0_n_50_16;
   wire execution_unit_0_n_50_17;
   wire execution_unit_0_n_50_18;
   wire execution_unit_0_n_50_19;
   wire execution_unit_0_n_50_20;
   wire execution_unit_0_n_50_21;
   wire execution_unit_0_n_50_22;
   wire execution_unit_0_n_50_23;
   wire execution_unit_0_n_50_24;
   wire execution_unit_0_n_50_25;
   wire execution_unit_0_n_50_26;
   wire execution_unit_0_n_50_27;
   wire execution_unit_0_n_50_28;
   wire execution_unit_0_n_50_29;
   wire execution_unit_0_n_50_30;
   wire execution_unit_0_n_50_31;
   wire execution_unit_0_n_50_32;
   wire execution_unit_0_n_50_33;
   wire execution_unit_0_n_50_34;
   wire execution_unit_0_n_50_35;
   wire execution_unit_0_n_50_36;
   wire execution_unit_0_n_50_37;
   wire execution_unit_0_n_50_38;
   wire execution_unit_0_n_50_39;
   wire execution_unit_0_n_50_40;
   wire execution_unit_0_n_50_41;
   wire execution_unit_0_n_50_42;
   wire execution_unit_0_n_50_43;
   wire execution_unit_0_n_50_44;
   wire execution_unit_0_n_50_45;
   wire execution_unit_0_n_50_46;
   wire execution_unit_0_n_50_47;
   wire execution_unit_0_n_50_48;
   wire execution_unit_0_n_50_49;
   wire execution_unit_0_n_50_50;
   wire execution_unit_0_n_50_51;
   wire execution_unit_0_n_50_52;
   wire execution_unit_0_n_50_53;
   wire execution_unit_0_n_50_54;
   wire execution_unit_0_n_50_55;
   wire execution_unit_0_n_50_56;
   wire execution_unit_0_n_50_57;
   wire execution_unit_0_n_50_58;
   wire execution_unit_0_n_50_59;
   wire execution_unit_0_n_50_60;
   wire execution_unit_0_n_50_61;
   wire execution_unit_0_n_50_62;
   wire execution_unit_0_n_50_63;
   wire execution_unit_0_n_50_64;
   wire execution_unit_0_n_50_65;
   wire execution_unit_0_n_50_66;
   wire execution_unit_0_n_50_67;
   wire execution_unit_0_n_50_68;
   wire execution_unit_0_n_50_69;
   wire execution_unit_0_n_50_70;
   wire execution_unit_0_n_50_71;
   wire execution_unit_0_n_50_72;
   wire execution_unit_0_n_50_73;
   wire execution_unit_0_n_50_74;
   wire execution_unit_0_n_50_75;
   wire execution_unit_0_n_50_76;
   wire execution_unit_0_n_50_77;
   wire execution_unit_0_n_50_78;
   wire execution_unit_0_n_50_79;
   wire execution_unit_0_n_50_80;
   wire execution_unit_0_n_50_81;
   wire execution_unit_0_n_50_82;
   wire execution_unit_0_n_50_83;
   wire execution_unit_0_n_50_84;
   wire execution_unit_0_n_50_85;
   wire execution_unit_0_n_50_86;
   wire execution_unit_0_n_50_87;
   wire execution_unit_0_n_50_88;
   wire execution_unit_0_n_50_89;
   wire execution_unit_0_n_50_90;
   wire execution_unit_0_n_50_91;
   wire execution_unit_0_n_50_92;
   wire execution_unit_0_n_50_93;
   wire execution_unit_0_n_50_94;
   wire execution_unit_0_n_50_95;
   wire execution_unit_0_n_0;
   wire execution_unit_0_n_69;
   wire execution_unit_0_n_1;
   wire execution_unit_0_n_2;
   wire execution_unit_0_n_73;
   wire execution_unit_0_n_74;
   wire execution_unit_0_n_3;
   wire execution_unit_0_n_40;
   wire execution_unit_0_n_10;
   wire execution_unit_0_n_67;
   wire execution_unit_0_n_68;
   wire execution_unit_0_n_72;
   wire execution_unit_0_n_75;
   wire execution_unit_0_n_47;
   wire execution_unit_0_n_13;
   wire execution_unit_0_n_11;
   wire execution_unit_0_n_6;
   wire execution_unit_0_n_5;
   wire execution_unit_0_n_12;
   wire execution_unit_0_n_4;
   wire execution_unit_0_n_9;
   wire execution_unit_0_n_16;
   wire execution_unit_0_n_18;
   wire execution_unit_0_n_49;
   wire execution_unit_0_n_48;
   wire execution_unit_0_n_65;
   wire execution_unit_0_n_37;
   wire execution_unit_0_n_38;
   wire execution_unit_0_n_71;
   wire execution_unit_0_n_76;
   wire execution_unit_0_n_41;
   wire execution_unit_0_n_42;
   wire execution_unit_0_n_43;
   wire execution_unit_0_n_8;
   wire execution_unit_0_n_44;
   wire execution_unit_0_n_46;
   wire execution_unit_0_n_66;
   wire execution_unit_0_n_7;
   wire execution_unit_0_n_45;
   wire execution_unit_0_n_70;
   wire execution_unit_0_n_77;
   wire execution_unit_0_n_93;
   wire execution_unit_0_n_64;
   wire execution_unit_0_n_92;
   wire execution_unit_0_n_63;
   wire execution_unit_0_n_91;
   wire execution_unit_0_n_62;
   wire execution_unit_0_n_90;
   wire execution_unit_0_n_61;
   wire execution_unit_0_n_89;
   wire execution_unit_0_n_60;
   wire execution_unit_0_n_88;
   wire execution_unit_0_n_59;
   wire execution_unit_0_n_87;
   wire execution_unit_0_n_58;
   wire execution_unit_0_n_86;
   wire execution_unit_0_n_57;
   wire execution_unit_0_n_85;
   wire execution_unit_0_n_56;
   wire execution_unit_0_n_84;
   wire execution_unit_0_n_55;
   wire execution_unit_0_n_83;
   wire execution_unit_0_n_54;
   wire execution_unit_0_n_82;
   wire execution_unit_0_n_53;
   wire execution_unit_0_n_81;
   wire execution_unit_0_n_52;
   wire execution_unit_0_n_80;
   wire execution_unit_0_n_51;
   wire execution_unit_0_n_79;
   wire execution_unit_0_n_50;
   wire execution_unit_0_n_78;
   wire execution_unit_0_n_102;
   wire execution_unit_0_n_98;
   wire execution_unit_0_n_103;
   wire execution_unit_0_n_96;
   wire execution_unit_0_n_97;
   wire execution_unit_0_n_95;
   wire execution_unit_0_n_101;
   wire execution_unit_0_n_105;
   wire execution_unit_0_n_94;
   wire execution_unit_0_n_106;
   wire execution_unit_0_n_39;
   wire execution_unit_0_n_100;
   wire execution_unit_0_n_107;
   wire execution_unit_0_n_99;
   wire execution_unit_0_n_108;
   wire execution_unit_0_n_104;
   wire execution_unit_0_n_124;
   wire execution_unit_0_n_123;
   wire execution_unit_0_n_122;
   wire execution_unit_0_n_121;
   wire execution_unit_0_n_120;
   wire execution_unit_0_n_119;
   wire execution_unit_0_n_118;
   wire execution_unit_0_n_117;
   wire execution_unit_0_n_116;
   wire execution_unit_0_n_115;
   wire execution_unit_0_n_114;
   wire execution_unit_0_n_113;
   wire execution_unit_0_n_112;
   wire execution_unit_0_n_111;
   wire execution_unit_0_n_110;
   wire execution_unit_0_n_109;
   wire execution_unit_0_n_15;
   wire execution_unit_0_n_14;
   wire execution_unit_0_n_34;
   wire execution_unit_0_n_35;
   wire execution_unit_0_n_36;
   wire execution_unit_0_n_17;
   wire execution_unit_0_n_26;
   wire execution_unit_0_n_33;
   wire execution_unit_0_n_25;
   wire execution_unit_0_n_32;
   wire execution_unit_0_n_24;
   wire execution_unit_0_n_31;
   wire execution_unit_0_n_23;
   wire execution_unit_0_n_30;
   wire execution_unit_0_n_22;
   wire execution_unit_0_n_29;
   wire execution_unit_0_n_21;
   wire execution_unit_0_n_28;
   wire execution_unit_0_n_20;
   wire execution_unit_0_n_27;
   wire execution_unit_0_n_19;
   wire execution_unit_0_alu_0_op_bit8_msk;
   wire execution_unit_0_alu_0_op_src_inv_cmd;
   wire execution_unit_0_alu_0_n_4_0;
   wire execution_unit_0_alu_0_n_4_1;
   wire execution_unit_0_alu_0_n_4_2;
   wire execution_unit_0_alu_0_n_4_3;
   wire execution_unit_0_alu_0_n_4_4;
   wire execution_unit_0_alu_0_n_4_5;
   wire [3:0]execution_unit_0_alu_0_X;
   wire execution_unit_0_alu_0_n_4_6;
   wire execution_unit_0_alu_0_n_4_7;
   wire execution_unit_0_alu_0_n_4_8;
   wire execution_unit_0_alu_0_n_5_0;
   wire execution_unit_0_alu_0_n_5_1;
   wire execution_unit_0_alu_0_n_5_2;
   wire execution_unit_0_alu_0_n_5_3;
   wire execution_unit_0_alu_0_n_5_4;
   wire execution_unit_0_alu_0_n_5_5;
   wire execution_unit_0_alu_0_n_6_0;
   wire execution_unit_0_alu_0_alu_short_thro;
   wire execution_unit_0_alu_0_n_7_0;
   wire execution_unit_0_alu_0_n_7_1;
   wire execution_unit_0_alu_0_n_7_2;
   wire execution_unit_0_alu_0_n_7_3;
   wire execution_unit_0_alu_0_n_7_4;
   wire execution_unit_0_alu_0_n_7_5;
   wire execution_unit_0_alu_0_n_7_6;
   wire execution_unit_0_alu_0_n_7_7;
   wire execution_unit_0_alu_0_n_7_8;
   wire execution_unit_0_alu_0_n_7_9;
   wire execution_unit_0_alu_0_n_7_10;
   wire execution_unit_0_alu_0_n_7_11;
   wire execution_unit_0_alu_0_n_7_12;
   wire execution_unit_0_alu_0_n_7_13;
   wire execution_unit_0_alu_0_n_7_14;
   wire execution_unit_0_alu_0_n_7_15;
   wire execution_unit_0_alu_0_n_7_16;
   wire execution_unit_0_alu_0_n_7_17;
   wire execution_unit_0_alu_0_n_7_18;
   wire execution_unit_0_alu_0_n_7_19;
   wire execution_unit_0_alu_0_n_7_20;
   wire execution_unit_0_alu_0_n_7_21;
   wire execution_unit_0_alu_0_n_7_22;
   wire execution_unit_0_alu_0_n_7_23;
   wire execution_unit_0_alu_0_n_7_24;
   wire execution_unit_0_alu_0_n_7_25;
   wire execution_unit_0_alu_0_n_7_26;
   wire execution_unit_0_alu_0_n_7_27;
   wire execution_unit_0_alu_0_n_7_28;
   wire execution_unit_0_alu_0_n_7_29;
   wire execution_unit_0_alu_0_n_7_30;
   wire execution_unit_0_alu_0_n_7_31;
   wire execution_unit_0_alu_0_n_7_32;
   wire execution_unit_0_alu_0_n_7_33;
   wire execution_unit_0_alu_0_n_7_34;
   wire execution_unit_0_alu_0_n_7_35;
   wire execution_unit_0_alu_0_n_7_36;
   wire execution_unit_0_alu_0_n_7_37;
   wire execution_unit_0_alu_0_n_7_38;
   wire execution_unit_0_alu_0_n_7_39;
   wire execution_unit_0_alu_0_n_7_40;
   wire execution_unit_0_alu_0_n_7_41;
   wire execution_unit_0_alu_0_n_7_42;
   wire execution_unit_0_alu_0_n_7_43;
   wire execution_unit_0_alu_0_n_7_44;
   wire execution_unit_0_alu_0_n_7_45;
   wire execution_unit_0_alu_0_n_7_46;
   wire execution_unit_0_alu_0_n_7_47;
   wire execution_unit_0_alu_0_n_7_48;
   wire execution_unit_0_alu_0_n_7_49;
   wire execution_unit_0_alu_0_n_7_50;
   wire execution_unit_0_alu_0_n_7_51;
   wire execution_unit_0_alu_0_n_7_52;
   wire execution_unit_0_alu_0_n_7_53;
   wire execution_unit_0_alu_0_n_7_54;
   wire execution_unit_0_alu_0_n_7_55;
   wire execution_unit_0_alu_0_n_7_56;
   wire execution_unit_0_alu_0_n_7_57;
   wire execution_unit_0_alu_0_n_7_58;
   wire execution_unit_0_alu_0_n_7_59;
   wire execution_unit_0_alu_0_n_7_60;
   wire execution_unit_0_alu_0_n_7_61;
   wire execution_unit_0_alu_0_n_7_62;
   wire execution_unit_0_alu_0_n_7_63;
   wire execution_unit_0_alu_0_n_7_64;
   wire execution_unit_0_alu_0_n_7_65;
   wire execution_unit_0_alu_0_n_7_66;
   wire execution_unit_0_alu_0_n_7_67;
   wire execution_unit_0_alu_0_n_7_68;
   wire execution_unit_0_alu_0_n_7_69;
   wire execution_unit_0_alu_0_n_7_70;
   wire execution_unit_0_alu_0_n_7_71;
   wire execution_unit_0_alu_0_n_7_72;
   wire execution_unit_0_alu_0_n_7_73;
   wire execution_unit_0_alu_0_n_7_74;
   wire execution_unit_0_alu_0_n_7_75;
   wire execution_unit_0_alu_0_n_7_76;
   wire execution_unit_0_alu_0_n_7_77;
   wire execution_unit_0_alu_0_n_7_78;
   wire execution_unit_0_alu_0_n_7_79;
   wire execution_unit_0_alu_0_n_7_80;
   wire execution_unit_0_alu_0_n_7_81;
   wire execution_unit_0_alu_0_n_7_82;
   wire execution_unit_0_alu_0_n_7_83;
   wire execution_unit_0_alu_0_n_7_84;
   wire execution_unit_0_alu_0_n_7_85;
   wire execution_unit_0_alu_0_n_7_86;
   wire execution_unit_0_alu_0_n_7_87;
   wire execution_unit_0_alu_0_n_7_88;
   wire execution_unit_0_alu_0_n_7_89;
   wire execution_unit_0_alu_0_n_7_90;
   wire execution_unit_0_alu_0_n_7_91;
   wire execution_unit_0_alu_0_n_7_92;
   wire execution_unit_0_alu_0_n_7_93;
   wire execution_unit_0_alu_0_n_7_94;
   wire execution_unit_0_alu_0_n_7_95;
   wire execution_unit_0_alu_0_n_7_96;
   wire execution_unit_0_alu_0_n_7_97;
   wire execution_unit_0_alu_0_n_7_98;
   wire execution_unit_0_alu_0_n_7_99;
   wire execution_unit_0_alu_0_n_7_100;
   wire execution_unit_0_alu_0_n_7_101;
   wire execution_unit_0_alu_0_n_7_102;
   wire execution_unit_0_alu_0_n_7_103;
   wire execution_unit_0_alu_0_n_7_104;
   wire execution_unit_0_alu_0_n_7_105;
   wire execution_unit_0_alu_0_n_7_106;
   wire execution_unit_0_alu_0_n_7_107;
   wire execution_unit_0_alu_0_n_7_108;
   wire execution_unit_0_alu_0_n_7_109;
   wire execution_unit_0_alu_0_n_7_110;
   wire execution_unit_0_alu_0_n_7_111;
   wire execution_unit_0_alu_0_n_7_112;
   wire execution_unit_0_alu_0_n_7_113;
   wire execution_unit_0_alu_0_n_7_114;
   wire execution_unit_0_alu_0_n_7_115;
   wire execution_unit_0_alu_0_n_7_116;
   wire execution_unit_0_alu_0_n_7_117;
   wire execution_unit_0_alu_0_n_7_118;
   wire execution_unit_0_alu_0_n_7_119;
   wire execution_unit_0_alu_0_n_7_120;
   wire execution_unit_0_alu_0_n_7_121;
   wire execution_unit_0_alu_0_n_7_122;
   wire execution_unit_0_alu_0_n_7_123;
   wire execution_unit_0_alu_0_n_7_124;
   wire execution_unit_0_alu_0_n_7_125;
   wire execution_unit_0_alu_0_n_7_126;
   wire execution_unit_0_alu_0_n_7_127;
   wire execution_unit_0_alu_0_n_7_128;
   wire execution_unit_0_alu_0_n_7_129;
   wire execution_unit_0_alu_0_n_7_130;
   wire execution_unit_0_alu_0_n_7_131;
   wire execution_unit_0_alu_0_n_7_132;
   wire execution_unit_0_alu_0_n_7_133;
   wire execution_unit_0_alu_0_n_7_134;
   wire execution_unit_0_alu_0_n_7_135;
   wire execution_unit_0_alu_0_n_8_0;
   wire execution_unit_0_alu_0_n_9_0;
   wire execution_unit_0_alu_0_n_9_1;
   wire execution_unit_0_alu_0_n_9_2;
   wire execution_unit_0_alu_0_n_9_3;
   wire execution_unit_0_alu_0_n_9_4;
   wire execution_unit_0_alu_0_n_9_5;
   wire execution_unit_0_alu_0_n_9_6;
   wire execution_unit_0_alu_0_n_9_7;
   wire execution_unit_0_alu_0_n_9_8;
   wire execution_unit_0_alu_0_n_9_9;
   wire execution_unit_0_alu_0_n_11_0;
   wire execution_unit_0_alu_0_n_11_1;
   wire execution_unit_0_alu_0_n_11_2;
   wire execution_unit_0_alu_0_n_12_0;
   wire [4:0]execution_unit_0_alu_0_bcd_add;
   wire execution_unit_0_alu_0_n_12_1;
   wire execution_unit_0_alu_0_n_12_2;
   wire execution_unit_0_alu_0_n_12_3;
   wire execution_unit_0_alu_0_n_12_4;
   wire execution_unit_0_alu_0_n_12_5;
   wire execution_unit_0_alu_0_n_12_6;
   wire execution_unit_0_alu_0_n_12_7;
   wire execution_unit_0_alu_0_n_12_8;
   wire execution_unit_0_alu_0_n_13_0;
   wire execution_unit_0_alu_0_n_14_0;
   wire execution_unit_0_alu_0_n_14_1;
   wire execution_unit_0_alu_0_n_14_2;
   wire execution_unit_0_alu_0_n_14_3;
   wire execution_unit_0_alu_0_n_14_4;
   wire execution_unit_0_alu_0_n_14_5;
   wire execution_unit_0_alu_0_n_14_6;
   wire execution_unit_0_alu_0_n_14_7;
   wire execution_unit_0_alu_0_n_14_8;
   wire execution_unit_0_alu_0_n_14_9;
   wire execution_unit_0_alu_0_n_16_0;
   wire execution_unit_0_alu_0_n_16_1;
   wire execution_unit_0_alu_0_n_16_2;
   wire execution_unit_0_alu_0_n_17_0;
   wire [4:0]execution_unit_0_alu_0_bcd_add0;
   wire execution_unit_0_alu_0_n_17_1;
   wire execution_unit_0_alu_0_n_17_2;
   wire execution_unit_0_alu_0_n_17_3;
   wire execution_unit_0_alu_0_n_17_4;
   wire execution_unit_0_alu_0_n_17_5;
   wire execution_unit_0_alu_0_n_17_6;
   wire execution_unit_0_alu_0_n_17_7;
   wire execution_unit_0_alu_0_n_17_8;
   wire execution_unit_0_alu_0_n_18_0;
   wire execution_unit_0_alu_0_n_19_0;
   wire execution_unit_0_alu_0_n_19_1;
   wire execution_unit_0_alu_0_n_19_2;
   wire execution_unit_0_alu_0_n_19_3;
   wire execution_unit_0_alu_0_n_19_4;
   wire execution_unit_0_alu_0_n_19_5;
   wire execution_unit_0_alu_0_n_19_6;
   wire execution_unit_0_alu_0_n_19_7;
   wire execution_unit_0_alu_0_n_19_8;
   wire execution_unit_0_alu_0_n_19_9;
   wire execution_unit_0_alu_0_n_21_0;
   wire execution_unit_0_alu_0_n_21_1;
   wire execution_unit_0_alu_0_n_21_2;
   wire execution_unit_0_alu_0_n_22_0;
   wire [4:0]execution_unit_0_alu_0_bcd_add1;
   wire execution_unit_0_alu_0_n_22_1;
   wire execution_unit_0_alu_0_n_22_2;
   wire execution_unit_0_alu_0_n_22_3;
   wire execution_unit_0_alu_0_n_22_4;
   wire execution_unit_0_alu_0_n_22_5;
   wire execution_unit_0_alu_0_n_22_6;
   wire execution_unit_0_alu_0_n_22_7;
   wire execution_unit_0_alu_0_n_22_8;
   wire execution_unit_0_alu_0_n_23_0;
   wire execution_unit_0_alu_0_n_24_0;
   wire execution_unit_0_alu_0_n_24_1;
   wire execution_unit_0_alu_0_n_24_2;
   wire execution_unit_0_alu_0_n_24_3;
   wire execution_unit_0_alu_0_n_24_4;
   wire execution_unit_0_alu_0_n_24_5;
   wire execution_unit_0_alu_0_n_24_6;
   wire execution_unit_0_alu_0_n_24_7;
   wire execution_unit_0_alu_0_n_24_8;
   wire execution_unit_0_alu_0_n_24_9;
   wire execution_unit_0_alu_0_n_26_0;
   wire execution_unit_0_alu_0_n_26_1;
   wire execution_unit_0_alu_0_n_26_2;
   wire execution_unit_0_alu_0_n_27_0;
   wire [4:0]execution_unit_0_alu_0_bcd_add2;
   wire execution_unit_0_alu_0_n_27_1;
   wire execution_unit_0_alu_0_n_27_2;
   wire execution_unit_0_alu_0_n_27_3;
   wire execution_unit_0_alu_0_n_27_4;
   wire execution_unit_0_alu_0_n_27_5;
   wire execution_unit_0_alu_0_n_27_6;
   wire execution_unit_0_alu_0_n_27_7;
   wire execution_unit_0_alu_0_n_27_8;
   wire execution_unit_0_alu_0_n_28_0;
   wire execution_unit_0_alu_0_n_28_1;
   wire execution_unit_0_alu_0_alu_inc;
   wire execution_unit_0_alu_0_n_30_0;
   wire execution_unit_0_alu_0_n_30_1;
   wire execution_unit_0_alu_0_n_30_2;
   wire execution_unit_0_alu_0_n_30_3;
   wire execution_unit_0_alu_0_n_30_4;
   wire execution_unit_0_alu_0_n_30_5;
   wire execution_unit_0_alu_0_n_30_6;
   wire execution_unit_0_alu_0_n_30_7;
   wire execution_unit_0_alu_0_n_30_8;
   wire execution_unit_0_alu_0_n_30_9;
   wire execution_unit_0_alu_0_n_40_0;
   wire execution_unit_0_alu_0_n_40_1;
   wire execution_unit_0_alu_0_n_40_2;
   wire execution_unit_0_alu_0_n_40_3;
   wire execution_unit_0_alu_0_n_40_4;
   wire execution_unit_0_alu_0_n_40_5;
   wire execution_unit_0_alu_0_n_40_6;
   wire execution_unit_0_alu_0_n_40_7;
   wire execution_unit_0_alu_0_n_40_8;
   wire execution_unit_0_alu_0_n_40_9;
   wire execution_unit_0_alu_0_n_40_10;
   wire execution_unit_0_alu_0_n_40_11;
   wire execution_unit_0_alu_0_n_40_12;
   wire execution_unit_0_alu_0_n_40_13;
   wire execution_unit_0_alu_0_n_40_14;
   wire [16:0]execution_unit_0_alu_0_alu_add;
   wire [16:0]execution_unit_0_alu_0_alu_add_inc;
   wire execution_unit_0_alu_0_n_41_0;
   wire execution_unit_0_alu_0_n_41_1;
   wire execution_unit_0_alu_0_n_41_2;
   wire execution_unit_0_alu_0_n_41_3;
   wire execution_unit_0_alu_0_n_41_4;
   wire execution_unit_0_alu_0_n_41_5;
   wire execution_unit_0_alu_0_n_41_6;
   wire execution_unit_0_alu_0_n_41_7;
   wire execution_unit_0_alu_0_n_41_8;
   wire execution_unit_0_alu_0_n_41_9;
   wire execution_unit_0_alu_0_n_41_10;
   wire execution_unit_0_alu_0_n_41_11;
   wire execution_unit_0_alu_0_n_41_12;
   wire execution_unit_0_alu_0_n_41_13;
   wire execution_unit_0_alu_0_n_41_14;
   wire execution_unit_0_alu_0_n_41_15;
   wire execution_unit_0_alu_0_n_41_16;
   wire execution_unit_0_alu_0_n_43_0;
   wire execution_unit_0_alu_0_n_44_0;
   wire execution_unit_0_alu_0_n_44_1;
   wire execution_unit_0_alu_0_n_44_2;
   wire execution_unit_0_alu_0_n_44_3;
   wire execution_unit_0_alu_0_n_44_4;
   wire execution_unit_0_alu_0_n_44_5;
   wire execution_unit_0_alu_0_n_44_6;
   wire execution_unit_0_alu_0_n_44_7;
   wire execution_unit_0_alu_0_n_44_8;
   wire execution_unit_0_alu_0_n_44_9;
   wire execution_unit_0_alu_0_n_44_10;
   wire execution_unit_0_alu_0_n_44_11;
   wire execution_unit_0_alu_0_n_44_12;
   wire execution_unit_0_alu_0_n_44_13;
   wire execution_unit_0_alu_0_n_44_14;
   wire execution_unit_0_alu_0_n_44_15;
   wire execution_unit_0_alu_0_n_44_16;
   wire execution_unit_0_alu_0_n_46_0;
   wire execution_unit_0_alu_0_n_46_1;
   wire execution_unit_0_alu_0_n_46_2;
   wire execution_unit_0_alu_0_n_48_0;
   wire execution_unit_0_alu_0_n_48_1;
   wire execution_unit_0_alu_0_n_48_2;
   wire execution_unit_0_alu_0_n_49_0;
   wire execution_unit_0_alu_0_n_49_1;
   wire execution_unit_0_alu_0_n_49_2;
   wire execution_unit_0_alu_0_n_49_3;
   wire execution_unit_0_alu_0_n_49_4;
   wire execution_unit_0_alu_0_n_49_5;
   wire execution_unit_0_alu_0_n_49_6;
   wire execution_unit_0_alu_0_n_49_7;
   wire execution_unit_0_alu_0_n_49_8;
   wire execution_unit_0_alu_0_n_49_9;
   wire execution_unit_0_alu_0_Z;
   wire execution_unit_0_alu_0_n_51_0;
   wire execution_unit_0_alu_0_n_51_1;
   wire execution_unit_0_alu_0_n_51_2;
   wire execution_unit_0_alu_0_n_51_3;
   wire execution_unit_0_alu_0_n_51_4;
   wire execution_unit_0_alu_0_n_51_5;
   wire execution_unit_0_alu_0_n_51_6;
   wire execution_unit_0_alu_0_n_51_7;
   wire execution_unit_0_alu_0_n_51_8;
   wire execution_unit_0_alu_0_n_51_9;
   wire execution_unit_0_alu_0_n_51_10;
   wire execution_unit_0_alu_0_n_51_11;
   wire execution_unit_0_alu_0_n_51_12;
   wire execution_unit_0_alu_0_n_51_13;
   wire execution_unit_0_alu_0_n_51_14;
   wire execution_unit_0_alu_0_n_51_15;
   wire execution_unit_0_alu_0_n_51_16;
   wire execution_unit_0_alu_0_n_51_17;
   wire execution_unit_0_alu_0_n_51_18;
   wire execution_unit_0_alu_0_n_51_19;
   wire execution_unit_0_alu_0_n_51_20;
   wire execution_unit_0_alu_0_n_51_21;
   wire execution_unit_0_alu_0_n_51_22;
   wire execution_unit_0_alu_0_n_104;
   wire execution_unit_0_alu_0_n_7;
   wire execution_unit_0_alu_0_n_86;
   wire execution_unit_0_alu_0_n_87;
   wire execution_unit_0_alu_0_n_103;
   wire execution_unit_0_alu_0_n_6;
   wire execution_unit_0_alu_0_n_102;
   wire execution_unit_0_alu_0_n_5;
   wire execution_unit_0_alu_0_n_101;
   wire execution_unit_0_alu_0_n_4;
   wire execution_unit_0_alu_0_n_100;
   wire execution_unit_0_alu_0_n_3;
   wire execution_unit_0_alu_0_n_19;
   wire execution_unit_0_alu_0_n_99;
   wire execution_unit_0_alu_0_n_2;
   wire execution_unit_0_alu_0_n_18;
   wire execution_unit_0_alu_0_n_98;
   wire execution_unit_0_alu_0_n_1;
   wire execution_unit_0_alu_0_n_17;
   wire execution_unit_0_alu_0_n_97;
   wire execution_unit_0_alu_0_n_0;
   wire execution_unit_0_alu_0_n_16;
   wire execution_unit_0_alu_0_n_96;
   wire execution_unit_0_alu_0_n_15;
   wire execution_unit_0_alu_0_n_95;
   wire execution_unit_0_alu_0_n_14;
   wire execution_unit_0_alu_0_n_94;
   wire execution_unit_0_alu_0_n_13;
   wire execution_unit_0_alu_0_n_93;
   wire execution_unit_0_alu_0_n_12;
   wire execution_unit_0_alu_0_n_92;
   wire execution_unit_0_alu_0_n_11;
   wire execution_unit_0_alu_0_n_91;
   wire execution_unit_0_alu_0_n_10;
   wire execution_unit_0_alu_0_n_90;
   wire execution_unit_0_alu_0_n_9;
   wire execution_unit_0_alu_0_n_89;
   wire execution_unit_0_alu_0_n_8;
   wire execution_unit_0_alu_0_n_88;
   wire execution_unit_0_alu_0_n_106;
   wire execution_unit_0_alu_0_n_68;
   wire execution_unit_0_alu_0_n_67;
   wire execution_unit_0_alu_0_n_66;
   wire execution_unit_0_alu_0_n_65;
   wire execution_unit_0_alu_0_n_56;
   wire execution_unit_0_alu_0_n_55;
   wire execution_unit_0_alu_0_n_54;
   wire execution_unit_0_alu_0_n_53;
   wire execution_unit_0_alu_0_n_44;
   wire execution_unit_0_alu_0_n_43;
   wire execution_unit_0_alu_0_n_42;
   wire execution_unit_0_alu_0_n_41;
   wire execution_unit_0_alu_0_n_38;
   wire execution_unit_0_alu_0_n_40;
   wire execution_unit_0_alu_0_n_39;
   wire execution_unit_0_alu_0_n_45;
   wire execution_unit_0_alu_0_n_46;
   wire execution_unit_0_alu_0_n_47;
   wire execution_unit_0_alu_0_n_48;
   wire execution_unit_0_alu_0_n_49;
   wire execution_unit_0_alu_0_n_50;
   wire execution_unit_0_alu_0_n_52;
   wire execution_unit_0_alu_0_n_51;
   wire execution_unit_0_alu_0_n_57;
   wire execution_unit_0_alu_0_n_58;
   wire execution_unit_0_alu_0_n_59;
   wire execution_unit_0_alu_0_n_60;
   wire execution_unit_0_alu_0_n_61;
   wire execution_unit_0_alu_0_n_62;
   wire execution_unit_0_alu_0_n_64;
   wire execution_unit_0_alu_0_n_63;
   wire execution_unit_0_alu_0_n_69;
   wire execution_unit_0_alu_0_n_70;
   wire execution_unit_0_alu_0_n_71;
   wire execution_unit_0_alu_0_n_72;
   wire execution_unit_0_alu_0_n_73;
   wire execution_unit_0_alu_0_n_74;
   wire execution_unit_0_alu_0_n_76;
   wire execution_unit_0_alu_0_n_75;
   wire execution_unit_0_alu_0_n_78;
   wire execution_unit_0_alu_0_n_77;
   wire execution_unit_0_alu_0_n_83;
   wire execution_unit_0_alu_0_n_80;
   wire execution_unit_0_alu_0_n_79;
   wire execution_unit_0_alu_0_n_81;
   wire execution_unit_0_alu_0_n_82;
   wire execution_unit_0_alu_0_n_84;
   wire execution_unit_0_alu_0_n_105;
   wire execution_unit_0_alu_0_n_20;
   wire execution_unit_0_alu_0_n_37;
   wire execution_unit_0_alu_0_n_36;
   wire execution_unit_0_alu_0_n_35;
   wire execution_unit_0_alu_0_n_34;
   wire execution_unit_0_alu_0_n_33;
   wire execution_unit_0_alu_0_n_32;
   wire execution_unit_0_alu_0_n_31;
   wire execution_unit_0_alu_0_n_30;
   wire execution_unit_0_alu_0_n_21;
   wire execution_unit_0_alu_0_n_29;
   wire execution_unit_0_alu_0_n_28;
   wire execution_unit_0_alu_0_n_27;
   wire execution_unit_0_alu_0_n_26;
   wire execution_unit_0_alu_0_n_25;
   wire execution_unit_0_alu_0_n_24;
   wire execution_unit_0_alu_0_n_23;
   wire execution_unit_0_alu_0_n_22;
   wire execution_unit_0_alu_0_n_108;
   wire execution_unit_0_alu_0_n_110;
   wire execution_unit_0_alu_0_n_109;
   wire execution_unit_0_alu_0_n_111;
   wire execution_unit_0_alu_0_n_112;
   wire execution_unit_0_alu_0_n_85;
   wire execution_unit_0_alu_0_n_107;
   wire execution_unit_0_register_file_0_n_0_0;
   wire execution_unit_0_register_file_0_n_1_0;
   wire execution_unit_0_register_file_0_r2_wr;
   wire execution_unit_0_register_file_0_n_2_0;
   wire execution_unit_0_register_file_0_n_2_1;
   wire [4:0]execution_unit_0_register_file_0_r2_nxt;
   wire execution_unit_0_register_file_0_n_2_2;
   wire execution_unit_0_register_file_0_n_2_3;
   wire execution_unit_0_register_file_0_n_2_4;
   wire execution_unit_0_register_file_0_n_5_0;
   wire execution_unit_0_register_file_0_n_5_1;
   wire execution_unit_0_register_file_0_n_5_2;
   wire execution_unit_0_register_file_0_n_5_3;
   wire execution_unit_0_register_file_0_n_5_4;
   wire execution_unit_0_register_file_0_n_5_5;
   wire execution_unit_0_register_file_0_n_5_6;
   wire execution_unit_0_register_file_0_n_5_7;
   wire execution_unit_0_register_file_0_n_5_8;
   wire execution_unit_0_register_file_0_n_5_9;
   wire execution_unit_0_register_file_0_n_5_10;
   wire execution_unit_0_register_file_0_n_5_11;
   wire execution_unit_0_register_file_0_n_5_12;
   wire execution_unit_0_register_file_0_n_5_13;
   wire execution_unit_0_register_file_0_n_5_14;
   wire execution_unit_0_register_file_0_n_5_15;
   wire execution_unit_0_register_file_0_n_5_16;
   wire execution_unit_0_register_file_0_n_6_0;
   wire execution_unit_0_register_file_0_n_8_0;
   wire execution_unit_0_register_file_0_n_9_0;
   wire execution_unit_0_register_file_0_n_10_0;
   wire execution_unit_0_register_file_0_inst_src_in;
   wire execution_unit_0_register_file_0_r1_inc;
   wire execution_unit_0_register_file_0_r1_wr;
   wire execution_unit_0_register_file_0_n_13_0;
   wire execution_unit_0_register_file_0_n_13_1;
   wire execution_unit_0_register_file_0_n_14_0;
   wire execution_unit_0_register_file_0_r3_wr;
   wire [15:0]execution_unit_0_register_file_0_r3;
   wire execution_unit_0_register_file_0_n_17_0;
   wire execution_unit_0_register_file_0_r4_inc;
   wire execution_unit_0_register_file_0_r4_wr;
   wire execution_unit_0_register_file_0_n_20_0;
   wire [15:0]execution_unit_0_register_file_0_reg_incr_val;
   wire execution_unit_0_register_file_0_n_22_0;
   wire execution_unit_0_register_file_0_n_22_1;
   wire execution_unit_0_register_file_0_n_22_2;
   wire execution_unit_0_register_file_0_n_22_3;
   wire execution_unit_0_register_file_0_n_22_4;
   wire execution_unit_0_register_file_0_n_22_5;
   wire execution_unit_0_register_file_0_n_22_6;
   wire execution_unit_0_register_file_0_n_22_7;
   wire execution_unit_0_register_file_0_n_22_8;
   wire execution_unit_0_register_file_0_n_22_9;
   wire execution_unit_0_register_file_0_n_22_10;
   wire execution_unit_0_register_file_0_n_22_11;
   wire execution_unit_0_register_file_0_n_22_12;
   wire execution_unit_0_register_file_0_n_22_13;
   wire execution_unit_0_register_file_0_n_22_14;
   wire execution_unit_0_register_file_0_n_22_15;
   wire [15:0]execution_unit_0_register_file_0_r4;
   wire execution_unit_0_register_file_0_n_24_0;
   wire execution_unit_0_register_file_0_n_24_1;
   wire execution_unit_0_register_file_0_n_24_2;
   wire execution_unit_0_register_file_0_n_24_3;
   wire execution_unit_0_register_file_0_n_24_4;
   wire execution_unit_0_register_file_0_n_24_5;
   wire execution_unit_0_register_file_0_n_24_6;
   wire execution_unit_0_register_file_0_n_24_7;
   wire execution_unit_0_register_file_0_n_24_8;
   wire execution_unit_0_register_file_0_n_24_9;
   wire execution_unit_0_register_file_0_n_24_10;
   wire execution_unit_0_register_file_0_n_24_11;
   wire execution_unit_0_register_file_0_n_24_12;
   wire execution_unit_0_register_file_0_n_24_13;
   wire execution_unit_0_register_file_0_n_24_14;
   wire execution_unit_0_register_file_0_n_24_15;
   wire execution_unit_0_register_file_0_n_24_16;
   wire execution_unit_0_register_file_0_n_25_0;
   wire execution_unit_0_register_file_0_n_25_1;
   wire execution_unit_0_register_file_0_n_27_0;
   wire execution_unit_0_register_file_0_r5_inc;
   wire execution_unit_0_register_file_0_r5_wr;
   wire [15:0]execution_unit_0_register_file_0_r5;
   wire execution_unit_0_register_file_0_n_31_0;
   wire execution_unit_0_register_file_0_n_31_1;
   wire execution_unit_0_register_file_0_n_31_2;
   wire execution_unit_0_register_file_0_n_31_3;
   wire execution_unit_0_register_file_0_n_31_4;
   wire execution_unit_0_register_file_0_n_31_5;
   wire execution_unit_0_register_file_0_n_31_6;
   wire execution_unit_0_register_file_0_n_31_7;
   wire execution_unit_0_register_file_0_n_31_8;
   wire execution_unit_0_register_file_0_n_31_9;
   wire execution_unit_0_register_file_0_n_31_10;
   wire execution_unit_0_register_file_0_n_31_11;
   wire execution_unit_0_register_file_0_n_31_12;
   wire execution_unit_0_register_file_0_n_31_13;
   wire execution_unit_0_register_file_0_n_31_14;
   wire execution_unit_0_register_file_0_n_31_15;
   wire execution_unit_0_register_file_0_n_31_16;
   wire execution_unit_0_register_file_0_n_32_0;
   wire execution_unit_0_register_file_0_n_32_1;
   wire execution_unit_0_register_file_0_n_34_0;
   wire execution_unit_0_register_file_0_r6_inc;
   wire execution_unit_0_register_file_0_r6_wr;
   wire [15:0]execution_unit_0_register_file_0_r6;
   wire execution_unit_0_register_file_0_n_38_0;
   wire execution_unit_0_register_file_0_n_38_1;
   wire execution_unit_0_register_file_0_n_38_2;
   wire execution_unit_0_register_file_0_n_38_3;
   wire execution_unit_0_register_file_0_n_38_4;
   wire execution_unit_0_register_file_0_n_38_5;
   wire execution_unit_0_register_file_0_n_38_6;
   wire execution_unit_0_register_file_0_n_38_7;
   wire execution_unit_0_register_file_0_n_38_8;
   wire execution_unit_0_register_file_0_n_38_9;
   wire execution_unit_0_register_file_0_n_38_10;
   wire execution_unit_0_register_file_0_n_38_11;
   wire execution_unit_0_register_file_0_n_38_12;
   wire execution_unit_0_register_file_0_n_38_13;
   wire execution_unit_0_register_file_0_n_38_14;
   wire execution_unit_0_register_file_0_n_38_15;
   wire execution_unit_0_register_file_0_n_38_16;
   wire execution_unit_0_register_file_0_n_39_0;
   wire execution_unit_0_register_file_0_n_39_1;
   wire execution_unit_0_register_file_0_n_41_0;
   wire execution_unit_0_register_file_0_r7_inc;
   wire execution_unit_0_register_file_0_r7_wr;
   wire [15:0]execution_unit_0_register_file_0_r7;
   wire execution_unit_0_register_file_0_n_45_0;
   wire execution_unit_0_register_file_0_n_45_1;
   wire execution_unit_0_register_file_0_n_45_2;
   wire execution_unit_0_register_file_0_n_45_3;
   wire execution_unit_0_register_file_0_n_45_4;
   wire execution_unit_0_register_file_0_n_45_5;
   wire execution_unit_0_register_file_0_n_45_6;
   wire execution_unit_0_register_file_0_n_45_7;
   wire execution_unit_0_register_file_0_n_45_8;
   wire execution_unit_0_register_file_0_n_45_9;
   wire execution_unit_0_register_file_0_n_45_10;
   wire execution_unit_0_register_file_0_n_45_11;
   wire execution_unit_0_register_file_0_n_45_12;
   wire execution_unit_0_register_file_0_n_45_13;
   wire execution_unit_0_register_file_0_n_45_14;
   wire execution_unit_0_register_file_0_n_45_15;
   wire execution_unit_0_register_file_0_n_45_16;
   wire execution_unit_0_register_file_0_n_46_0;
   wire execution_unit_0_register_file_0_n_46_1;
   wire execution_unit_0_register_file_0_n_48_0;
   wire execution_unit_0_register_file_0_r8_inc;
   wire execution_unit_0_register_file_0_r8_wr;
   wire [15:0]execution_unit_0_register_file_0_r8;
   wire execution_unit_0_register_file_0_n_52_0;
   wire execution_unit_0_register_file_0_n_52_1;
   wire execution_unit_0_register_file_0_n_52_2;
   wire execution_unit_0_register_file_0_n_52_3;
   wire execution_unit_0_register_file_0_n_52_4;
   wire execution_unit_0_register_file_0_n_52_5;
   wire execution_unit_0_register_file_0_n_52_6;
   wire execution_unit_0_register_file_0_n_52_7;
   wire execution_unit_0_register_file_0_n_52_8;
   wire execution_unit_0_register_file_0_n_52_9;
   wire execution_unit_0_register_file_0_n_52_10;
   wire execution_unit_0_register_file_0_n_52_11;
   wire execution_unit_0_register_file_0_n_52_12;
   wire execution_unit_0_register_file_0_n_52_13;
   wire execution_unit_0_register_file_0_n_52_14;
   wire execution_unit_0_register_file_0_n_52_15;
   wire execution_unit_0_register_file_0_n_52_16;
   wire execution_unit_0_register_file_0_n_53_0;
   wire execution_unit_0_register_file_0_n_53_1;
   wire execution_unit_0_register_file_0_n_55_0;
   wire execution_unit_0_register_file_0_r9_inc;
   wire execution_unit_0_register_file_0_r9_wr;
   wire [15:0]execution_unit_0_register_file_0_r9;
   wire execution_unit_0_register_file_0_n_59_0;
   wire execution_unit_0_register_file_0_n_59_1;
   wire execution_unit_0_register_file_0_n_59_2;
   wire execution_unit_0_register_file_0_n_59_3;
   wire execution_unit_0_register_file_0_n_59_4;
   wire execution_unit_0_register_file_0_n_59_5;
   wire execution_unit_0_register_file_0_n_59_6;
   wire execution_unit_0_register_file_0_n_59_7;
   wire execution_unit_0_register_file_0_n_59_8;
   wire execution_unit_0_register_file_0_n_59_9;
   wire execution_unit_0_register_file_0_n_59_10;
   wire execution_unit_0_register_file_0_n_59_11;
   wire execution_unit_0_register_file_0_n_59_12;
   wire execution_unit_0_register_file_0_n_59_13;
   wire execution_unit_0_register_file_0_n_59_14;
   wire execution_unit_0_register_file_0_n_59_15;
   wire execution_unit_0_register_file_0_n_59_16;
   wire execution_unit_0_register_file_0_n_60_0;
   wire execution_unit_0_register_file_0_n_60_1;
   wire execution_unit_0_register_file_0_n_62_0;
   wire execution_unit_0_register_file_0_r10_inc;
   wire execution_unit_0_register_file_0_r10_wr;
   wire [15:0]execution_unit_0_register_file_0_r10;
   wire execution_unit_0_register_file_0_n_66_0;
   wire execution_unit_0_register_file_0_n_66_1;
   wire execution_unit_0_register_file_0_n_66_2;
   wire execution_unit_0_register_file_0_n_66_3;
   wire execution_unit_0_register_file_0_n_66_4;
   wire execution_unit_0_register_file_0_n_66_5;
   wire execution_unit_0_register_file_0_n_66_6;
   wire execution_unit_0_register_file_0_n_66_7;
   wire execution_unit_0_register_file_0_n_66_8;
   wire execution_unit_0_register_file_0_n_66_9;
   wire execution_unit_0_register_file_0_n_66_10;
   wire execution_unit_0_register_file_0_n_66_11;
   wire execution_unit_0_register_file_0_n_66_12;
   wire execution_unit_0_register_file_0_n_66_13;
   wire execution_unit_0_register_file_0_n_66_14;
   wire execution_unit_0_register_file_0_n_66_15;
   wire execution_unit_0_register_file_0_n_66_16;
   wire execution_unit_0_register_file_0_n_67_0;
   wire execution_unit_0_register_file_0_n_67_1;
   wire execution_unit_0_register_file_0_n_69_0;
   wire execution_unit_0_register_file_0_r11_inc;
   wire execution_unit_0_register_file_0_r11_wr;
   wire [15:0]execution_unit_0_register_file_0_r11;
   wire execution_unit_0_register_file_0_n_73_0;
   wire execution_unit_0_register_file_0_n_73_1;
   wire execution_unit_0_register_file_0_n_73_2;
   wire execution_unit_0_register_file_0_n_73_3;
   wire execution_unit_0_register_file_0_n_73_4;
   wire execution_unit_0_register_file_0_n_73_5;
   wire execution_unit_0_register_file_0_n_73_6;
   wire execution_unit_0_register_file_0_n_73_7;
   wire execution_unit_0_register_file_0_n_73_8;
   wire execution_unit_0_register_file_0_n_73_9;
   wire execution_unit_0_register_file_0_n_73_10;
   wire execution_unit_0_register_file_0_n_73_11;
   wire execution_unit_0_register_file_0_n_73_12;
   wire execution_unit_0_register_file_0_n_73_13;
   wire execution_unit_0_register_file_0_n_73_14;
   wire execution_unit_0_register_file_0_n_73_15;
   wire execution_unit_0_register_file_0_n_73_16;
   wire execution_unit_0_register_file_0_n_74_0;
   wire execution_unit_0_register_file_0_n_74_1;
   wire execution_unit_0_register_file_0_n_76_0;
   wire execution_unit_0_register_file_0_r12_inc;
   wire execution_unit_0_register_file_0_r12_wr;
   wire [15:0]execution_unit_0_register_file_0_r12;
   wire execution_unit_0_register_file_0_n_80_0;
   wire execution_unit_0_register_file_0_n_80_1;
   wire execution_unit_0_register_file_0_n_80_2;
   wire execution_unit_0_register_file_0_n_80_3;
   wire execution_unit_0_register_file_0_n_80_4;
   wire execution_unit_0_register_file_0_n_80_5;
   wire execution_unit_0_register_file_0_n_80_6;
   wire execution_unit_0_register_file_0_n_80_7;
   wire execution_unit_0_register_file_0_n_80_8;
   wire execution_unit_0_register_file_0_n_80_9;
   wire execution_unit_0_register_file_0_n_80_10;
   wire execution_unit_0_register_file_0_n_80_11;
   wire execution_unit_0_register_file_0_n_80_12;
   wire execution_unit_0_register_file_0_n_80_13;
   wire execution_unit_0_register_file_0_n_80_14;
   wire execution_unit_0_register_file_0_n_80_15;
   wire execution_unit_0_register_file_0_n_80_16;
   wire execution_unit_0_register_file_0_n_81_0;
   wire execution_unit_0_register_file_0_n_81_1;
   wire execution_unit_0_register_file_0_n_83_0;
   wire execution_unit_0_register_file_0_r13_inc;
   wire execution_unit_0_register_file_0_r13_wr;
   wire [15:0]execution_unit_0_register_file_0_r13;
   wire execution_unit_0_register_file_0_n_87_0;
   wire execution_unit_0_register_file_0_n_87_1;
   wire execution_unit_0_register_file_0_n_87_2;
   wire execution_unit_0_register_file_0_n_87_3;
   wire execution_unit_0_register_file_0_n_87_4;
   wire execution_unit_0_register_file_0_n_87_5;
   wire execution_unit_0_register_file_0_n_87_6;
   wire execution_unit_0_register_file_0_n_87_7;
   wire execution_unit_0_register_file_0_n_87_8;
   wire execution_unit_0_register_file_0_n_87_9;
   wire execution_unit_0_register_file_0_n_87_10;
   wire execution_unit_0_register_file_0_n_87_11;
   wire execution_unit_0_register_file_0_n_87_12;
   wire execution_unit_0_register_file_0_n_87_13;
   wire execution_unit_0_register_file_0_n_87_14;
   wire execution_unit_0_register_file_0_n_87_15;
   wire execution_unit_0_register_file_0_n_87_16;
   wire execution_unit_0_register_file_0_n_88_0;
   wire execution_unit_0_register_file_0_n_88_1;
   wire execution_unit_0_register_file_0_n_90_0;
   wire execution_unit_0_register_file_0_r14_inc;
   wire execution_unit_0_register_file_0_r14_wr;
   wire [15:0]execution_unit_0_register_file_0_r14;
   wire execution_unit_0_register_file_0_n_94_0;
   wire execution_unit_0_register_file_0_n_94_1;
   wire execution_unit_0_register_file_0_n_94_2;
   wire execution_unit_0_register_file_0_n_94_3;
   wire execution_unit_0_register_file_0_n_94_4;
   wire execution_unit_0_register_file_0_n_94_5;
   wire execution_unit_0_register_file_0_n_94_6;
   wire execution_unit_0_register_file_0_n_94_7;
   wire execution_unit_0_register_file_0_n_94_8;
   wire execution_unit_0_register_file_0_n_94_9;
   wire execution_unit_0_register_file_0_n_94_10;
   wire execution_unit_0_register_file_0_n_94_11;
   wire execution_unit_0_register_file_0_n_94_12;
   wire execution_unit_0_register_file_0_n_94_13;
   wire execution_unit_0_register_file_0_n_94_14;
   wire execution_unit_0_register_file_0_n_94_15;
   wire execution_unit_0_register_file_0_n_94_16;
   wire execution_unit_0_register_file_0_n_95_0;
   wire execution_unit_0_register_file_0_n_95_1;
   wire execution_unit_0_register_file_0_n_97_0;
   wire execution_unit_0_register_file_0_r15_inc;
   wire execution_unit_0_register_file_0_r15_wr;
   wire [15:0]execution_unit_0_register_file_0_r15;
   wire execution_unit_0_register_file_0_n_101_0;
   wire execution_unit_0_register_file_0_n_101_1;
   wire execution_unit_0_register_file_0_n_101_2;
   wire execution_unit_0_register_file_0_n_101_3;
   wire execution_unit_0_register_file_0_n_101_4;
   wire execution_unit_0_register_file_0_n_101_5;
   wire execution_unit_0_register_file_0_n_101_6;
   wire execution_unit_0_register_file_0_n_101_7;
   wire execution_unit_0_register_file_0_n_101_8;
   wire execution_unit_0_register_file_0_n_101_9;
   wire execution_unit_0_register_file_0_n_101_10;
   wire execution_unit_0_register_file_0_n_101_11;
   wire execution_unit_0_register_file_0_n_101_12;
   wire execution_unit_0_register_file_0_n_101_13;
   wire execution_unit_0_register_file_0_n_101_14;
   wire execution_unit_0_register_file_0_n_101_15;
   wire execution_unit_0_register_file_0_n_101_16;
   wire execution_unit_0_register_file_0_n_102_0;
   wire execution_unit_0_register_file_0_n_102_1;
   wire execution_unit_0_register_file_0_n_104_0;
   wire execution_unit_0_register_file_0_n_105_0;
   wire execution_unit_0_register_file_0_n_105_1;
   wire execution_unit_0_register_file_0_n_105_2;
   wire execution_unit_0_register_file_0_n_105_3;
   wire execution_unit_0_register_file_0_n_105_4;
   wire execution_unit_0_register_file_0_n_105_5;
   wire execution_unit_0_register_file_0_n_105_6;
   wire execution_unit_0_register_file_0_n_105_7;
   wire execution_unit_0_register_file_0_n_105_8;
   wire execution_unit_0_register_file_0_n_105_9;
   wire execution_unit_0_register_file_0_n_105_10;
   wire execution_unit_0_register_file_0_n_105_11;
   wire execution_unit_0_register_file_0_n_105_12;
   wire execution_unit_0_register_file_0_n_105_13;
   wire execution_unit_0_register_file_0_n_105_14;
   wire execution_unit_0_register_file_0_n_105_15;
   wire execution_unit_0_register_file_0_n_105_16;
   wire execution_unit_0_register_file_0_n_105_17;
   wire execution_unit_0_register_file_0_n_105_18;
   wire execution_unit_0_register_file_0_n_105_19;
   wire execution_unit_0_register_file_0_n_105_20;
   wire execution_unit_0_register_file_0_n_105_21;
   wire execution_unit_0_register_file_0_n_105_22;
   wire execution_unit_0_register_file_0_n_105_23;
   wire execution_unit_0_register_file_0_n_105_24;
   wire execution_unit_0_register_file_0_n_105_25;
   wire execution_unit_0_register_file_0_n_105_26;
   wire execution_unit_0_register_file_0_n_105_27;
   wire execution_unit_0_register_file_0_n_105_28;
   wire execution_unit_0_register_file_0_n_105_29;
   wire execution_unit_0_register_file_0_n_105_30;
   wire execution_unit_0_register_file_0_n_105_31;
   wire execution_unit_0_register_file_0_n_105_32;
   wire execution_unit_0_register_file_0_n_105_33;
   wire execution_unit_0_register_file_0_n_105_34;
   wire execution_unit_0_register_file_0_n_105_35;
   wire execution_unit_0_register_file_0_n_105_36;
   wire execution_unit_0_register_file_0_n_105_37;
   wire execution_unit_0_register_file_0_n_105_38;
   wire execution_unit_0_register_file_0_n_105_39;
   wire execution_unit_0_register_file_0_n_105_40;
   wire execution_unit_0_register_file_0_n_105_41;
   wire execution_unit_0_register_file_0_n_105_42;
   wire execution_unit_0_register_file_0_n_105_43;
   wire execution_unit_0_register_file_0_n_105_44;
   wire execution_unit_0_register_file_0_n_105_45;
   wire execution_unit_0_register_file_0_n_105_46;
   wire execution_unit_0_register_file_0_n_105_47;
   wire execution_unit_0_register_file_0_n_105_48;
   wire execution_unit_0_register_file_0_n_105_49;
   wire execution_unit_0_register_file_0_n_105_50;
   wire execution_unit_0_register_file_0_n_105_51;
   wire execution_unit_0_register_file_0_n_105_52;
   wire execution_unit_0_register_file_0_n_105_53;
   wire execution_unit_0_register_file_0_n_105_54;
   wire execution_unit_0_register_file_0_n_105_55;
   wire execution_unit_0_register_file_0_n_105_56;
   wire execution_unit_0_register_file_0_n_105_57;
   wire execution_unit_0_register_file_0_n_105_58;
   wire execution_unit_0_register_file_0_n_105_59;
   wire execution_unit_0_register_file_0_n_105_60;
   wire execution_unit_0_register_file_0_n_105_61;
   wire execution_unit_0_register_file_0_n_105_62;
   wire execution_unit_0_register_file_0_n_105_63;
   wire execution_unit_0_register_file_0_n_105_64;
   wire execution_unit_0_register_file_0_n_105_65;
   wire execution_unit_0_register_file_0_n_105_66;
   wire execution_unit_0_register_file_0_n_105_67;
   wire execution_unit_0_register_file_0_n_105_68;
   wire execution_unit_0_register_file_0_n_105_69;
   wire execution_unit_0_register_file_0_n_105_70;
   wire execution_unit_0_register_file_0_n_105_71;
   wire execution_unit_0_register_file_0_n_105_72;
   wire execution_unit_0_register_file_0_n_105_73;
   wire execution_unit_0_register_file_0_n_105_74;
   wire execution_unit_0_register_file_0_n_105_75;
   wire execution_unit_0_register_file_0_n_105_76;
   wire execution_unit_0_register_file_0_n_105_77;
   wire execution_unit_0_register_file_0_n_105_78;
   wire execution_unit_0_register_file_0_n_105_79;
   wire execution_unit_0_register_file_0_n_105_80;
   wire execution_unit_0_register_file_0_n_105_81;
   wire execution_unit_0_register_file_0_n_105_82;
   wire execution_unit_0_register_file_0_n_105_83;
   wire execution_unit_0_register_file_0_n_105_84;
   wire execution_unit_0_register_file_0_n_105_85;
   wire execution_unit_0_register_file_0_n_105_86;
   wire execution_unit_0_register_file_0_n_105_87;
   wire execution_unit_0_register_file_0_n_105_88;
   wire execution_unit_0_register_file_0_n_105_89;
   wire execution_unit_0_register_file_0_n_105_90;
   wire execution_unit_0_register_file_0_n_105_91;
   wire execution_unit_0_register_file_0_n_105_92;
   wire execution_unit_0_register_file_0_n_105_93;
   wire execution_unit_0_register_file_0_n_105_94;
   wire execution_unit_0_register_file_0_n_105_95;
   wire execution_unit_0_register_file_0_n_105_96;
   wire execution_unit_0_register_file_0_n_105_97;
   wire execution_unit_0_register_file_0_n_105_98;
   wire execution_unit_0_register_file_0_n_105_99;
   wire execution_unit_0_register_file_0_n_105_100;
   wire execution_unit_0_register_file_0_n_105_101;
   wire execution_unit_0_register_file_0_n_105_102;
   wire execution_unit_0_register_file_0_n_105_103;
   wire execution_unit_0_register_file_0_n_105_104;
   wire execution_unit_0_register_file_0_n_105_105;
   wire execution_unit_0_register_file_0_n_105_106;
   wire execution_unit_0_register_file_0_n_105_107;
   wire execution_unit_0_register_file_0_n_105_108;
   wire execution_unit_0_register_file_0_n_105_109;
   wire execution_unit_0_register_file_0_n_105_110;
   wire execution_unit_0_register_file_0_n_105_111;
   wire execution_unit_0_register_file_0_n_105_112;
   wire execution_unit_0_register_file_0_n_105_113;
   wire execution_unit_0_register_file_0_n_105_114;
   wire execution_unit_0_register_file_0_n_105_115;
   wire execution_unit_0_register_file_0_n_105_116;
   wire execution_unit_0_register_file_0_n_105_117;
   wire execution_unit_0_register_file_0_n_105_118;
   wire execution_unit_0_register_file_0_n_105_119;
   wire execution_unit_0_register_file_0_n_105_120;
   wire execution_unit_0_register_file_0_n_105_121;
   wire execution_unit_0_register_file_0_n_105_122;
   wire execution_unit_0_register_file_0_n_105_123;
   wire execution_unit_0_register_file_0_n_105_124;
   wire execution_unit_0_register_file_0_n_105_125;
   wire execution_unit_0_register_file_0_n_105_126;
   wire execution_unit_0_register_file_0_n_105_127;
   wire execution_unit_0_register_file_0_n_105_128;
   wire execution_unit_0_register_file_0_n_105_129;
   wire execution_unit_0_register_file_0_n_105_130;
   wire execution_unit_0_register_file_0_n_105_131;
   wire execution_unit_0_register_file_0_n_105_132;
   wire execution_unit_0_register_file_0_n_105_133;
   wire execution_unit_0_register_file_0_n_105_134;
   wire execution_unit_0_register_file_0_n_105_135;
   wire execution_unit_0_register_file_0_n_105_136;
   wire execution_unit_0_register_file_0_n_105_137;
   wire execution_unit_0_register_file_0_n_105_138;
   wire execution_unit_0_register_file_0_n_105_139;
   wire execution_unit_0_register_file_0_n_105_140;
   wire execution_unit_0_register_file_0_n_105_141;
   wire execution_unit_0_register_file_0_n_105_142;
   wire execution_unit_0_register_file_0_n_105_143;
   wire execution_unit_0_register_file_0_n_105_144;
   wire execution_unit_0_register_file_0_n_105_145;
   wire execution_unit_0_register_file_0_n_105_146;
   wire execution_unit_0_register_file_0_n_105_147;
   wire execution_unit_0_register_file_0_n_105_148;
   wire execution_unit_0_register_file_0_n_105_149;
   wire execution_unit_0_register_file_0_n_105_150;
   wire execution_unit_0_register_file_0_n_105_151;
   wire execution_unit_0_register_file_0_n_105_152;
   wire execution_unit_0_register_file_0_n_105_153;
   wire execution_unit_0_register_file_0_n_105_154;
   wire execution_unit_0_register_file_0_n_105_155;
   wire execution_unit_0_register_file_0_n_105_156;
   wire execution_unit_0_register_file_0_n_105_157;
   wire execution_unit_0_register_file_0_n_105_158;
   wire execution_unit_0_register_file_0_n_105_159;
   wire execution_unit_0_register_file_0_n_105_160;
   wire execution_unit_0_register_file_0_n_105_161;
   wire execution_unit_0_register_file_0_n_105_162;
   wire execution_unit_0_register_file_0_n_105_163;
   wire execution_unit_0_register_file_0_n_105_164;
   wire execution_unit_0_register_file_0_n_105_165;
   wire execution_unit_0_register_file_0_n_105_166;
   wire execution_unit_0_register_file_0_n_105_167;
   wire execution_unit_0_register_file_0_n_105_168;
   wire execution_unit_0_register_file_0_n_105_169;
   wire execution_unit_0_register_file_0_n_105_170;
   wire execution_unit_0_register_file_0_n_105_171;
   wire execution_unit_0_register_file_0_n_105_172;
   wire execution_unit_0_register_file_0_n_105_173;
   wire execution_unit_0_register_file_0_n_105_174;
   wire execution_unit_0_register_file_0_n_105_175;
   wire execution_unit_0_register_file_0_n_105_176;
   wire execution_unit_0_register_file_0_n_105_177;
   wire execution_unit_0_register_file_0_n_105_178;
   wire execution_unit_0_register_file_0_n_105_179;
   wire execution_unit_0_register_file_0_n_105_180;
   wire execution_unit_0_register_file_0_n_105_181;
   wire execution_unit_0_register_file_0_n_105_182;
   wire execution_unit_0_register_file_0_n_105_183;
   wire execution_unit_0_register_file_0_n_105_184;
   wire execution_unit_0_register_file_0_n_105_185;
   wire execution_unit_0_register_file_0_n_105_186;
   wire execution_unit_0_register_file_0_n_105_187;
   wire execution_unit_0_register_file_0_n_105_188;
   wire execution_unit_0_register_file_0_n_105_189;
   wire execution_unit_0_register_file_0_n_105_190;
   wire execution_unit_0_register_file_0_n_105_191;
   wire execution_unit_0_register_file_0_n_105_192;
   wire execution_unit_0_register_file_0_n_105_193;
   wire execution_unit_0_register_file_0_n_105_194;
   wire execution_unit_0_register_file_0_n_105_195;
   wire execution_unit_0_register_file_0_n_105_196;
   wire execution_unit_0_register_file_0_n_105_197;
   wire execution_unit_0_register_file_0_n_105_198;
   wire execution_unit_0_register_file_0_n_105_199;
   wire execution_unit_0_register_file_0_n_105_200;
   wire execution_unit_0_register_file_0_n_105_201;
   wire execution_unit_0_register_file_0_n_105_202;
   wire execution_unit_0_register_file_0_n_105_203;
   wire execution_unit_0_register_file_0_n_105_204;
   wire execution_unit_0_register_file_0_n_105_205;
   wire execution_unit_0_register_file_0_n_105_206;
   wire execution_unit_0_register_file_0_n_105_207;
   wire execution_unit_0_register_file_0_n_105_208;
   wire execution_unit_0_register_file_0_n_105_209;
   wire execution_unit_0_register_file_0_n_105_210;
   wire execution_unit_0_register_file_0_n_105_211;
   wire execution_unit_0_register_file_0_n_105_212;
   wire execution_unit_0_register_file_0_n_105_213;
   wire execution_unit_0_register_file_0_n_105_214;
   wire execution_unit_0_register_file_0_n_105_215;
   wire execution_unit_0_register_file_0_n_105_216;
   wire execution_unit_0_register_file_0_n_105_217;
   wire execution_unit_0_register_file_0_n_105_218;
   wire execution_unit_0_register_file_0_n_105_219;
   wire execution_unit_0_register_file_0_n_105_220;
   wire execution_unit_0_register_file_0_n_105_221;
   wire execution_unit_0_register_file_0_n_105_222;
   wire execution_unit_0_register_file_0_n_105_223;
   wire execution_unit_0_register_file_0_n_105_224;
   wire execution_unit_0_register_file_0_n_105_225;
   wire execution_unit_0_register_file_0_n_105_226;
   wire execution_unit_0_register_file_0_n_105_227;
   wire execution_unit_0_register_file_0_n_105_228;
   wire execution_unit_0_register_file_0_n_105_229;
   wire execution_unit_0_register_file_0_n_105_230;
   wire execution_unit_0_register_file_0_n_105_231;
   wire execution_unit_0_register_file_0_n_105_232;
   wire execution_unit_0_register_file_0_n_105_233;
   wire execution_unit_0_register_file_0_n_105_234;
   wire execution_unit_0_register_file_0_n_105_235;
   wire execution_unit_0_register_file_0_n_105_236;
   wire execution_unit_0_register_file_0_n_105_237;
   wire execution_unit_0_register_file_0_n_105_238;
   wire execution_unit_0_register_file_0_n_105_239;
   wire execution_unit_0_register_file_0_n_105_240;
   wire execution_unit_0_register_file_0_n_105_241;
   wire execution_unit_0_register_file_0_n_105_242;
   wire execution_unit_0_register_file_0_n_105_243;
   wire execution_unit_0_register_file_0_n_105_244;
   wire execution_unit_0_register_file_0_n_105_245;
   wire execution_unit_0_register_file_0_n_105_246;
   wire execution_unit_0_register_file_0_n_105_247;
   wire execution_unit_0_register_file_0_n_105_248;
   wire execution_unit_0_register_file_0_n_105_249;
   wire execution_unit_0_register_file_0_n_105_250;
   wire execution_unit_0_register_file_0_n_105_251;
   wire execution_unit_0_register_file_0_n_105_252;
   wire execution_unit_0_register_file_0_n_105_253;
   wire execution_unit_0_register_file_0_n_105_254;
   wire execution_unit_0_register_file_0_n_105_255;
   wire execution_unit_0_register_file_0_n_105_256;
   wire execution_unit_0_register_file_0_n_105_257;
   wire execution_unit_0_register_file_0_n_105_258;
   wire execution_unit_0_register_file_0_n_105_259;
   wire execution_unit_0_register_file_0_n_105_260;
   wire execution_unit_0_register_file_0_n_105_261;
   wire execution_unit_0_register_file_0_n_105_262;
   wire execution_unit_0_register_file_0_n_105_263;
   wire execution_unit_0_register_file_0_n_105_264;
   wire execution_unit_0_register_file_0_n_105_265;
   wire execution_unit_0_register_file_0_n_105_266;
   wire execution_unit_0_register_file_0_n_105_267;
   wire execution_unit_0_register_file_0_n_105_268;
   wire execution_unit_0_register_file_0_n_105_269;
   wire execution_unit_0_register_file_0_n_105_270;
   wire execution_unit_0_register_file_0_n_105_271;
   wire execution_unit_0_register_file_0_n_105_272;
   wire execution_unit_0_register_file_0_n_105_273;
   wire execution_unit_0_register_file_0_n_105_274;
   wire execution_unit_0_register_file_0_n_105_275;
   wire execution_unit_0_register_file_0_n_105_276;
   wire execution_unit_0_register_file_0_n_105_277;
   wire execution_unit_0_register_file_0_n_105_278;
   wire execution_unit_0_register_file_0_n_105_279;
   wire execution_unit_0_register_file_0_n_105_280;
   wire execution_unit_0_register_file_0_n_105_281;
   wire execution_unit_0_register_file_0_n_105_282;
   wire execution_unit_0_register_file_0_n_105_283;
   wire execution_unit_0_register_file_0_n_105_284;
   wire execution_unit_0_register_file_0_n_105_285;
   wire execution_unit_0_register_file_0_n_105_286;
   wire execution_unit_0_register_file_0_n_105_287;
   wire execution_unit_0_register_file_0_n_105_288;
   wire execution_unit_0_register_file_0_n_105_289;
   wire execution_unit_0_register_file_0_n_105_290;
   wire execution_unit_0_register_file_0_n_105_291;
   wire execution_unit_0_register_file_0_n_105_292;
   wire execution_unit_0_register_file_0_n_105_293;
   wire execution_unit_0_register_file_0_n_105_294;
   wire execution_unit_0_register_file_0_n_105_295;
   wire execution_unit_0_register_file_0_n_105_296;
   wire execution_unit_0_register_file_0_n_105_297;
   wire execution_unit_0_register_file_0_n_105_298;
   wire execution_unit_0_register_file_0_n_105_299;
   wire execution_unit_0_register_file_0_n_105_300;
   wire execution_unit_0_register_file_0_n_105_301;
   wire execution_unit_0_register_file_0_n_105_302;
   wire execution_unit_0_register_file_0_n_105_303;
   wire execution_unit_0_register_file_0_n_105_304;
   wire execution_unit_0_register_file_0_n_105_305;
   wire execution_unit_0_register_file_0_n_105_306;
   wire execution_unit_0_register_file_0_n_105_307;
   wire execution_unit_0_register_file_0_n_105_308;
   wire execution_unit_0_register_file_0_n_105_309;
   wire execution_unit_0_register_file_0_n_105_310;
   wire execution_unit_0_register_file_0_n_105_311;
   wire execution_unit_0_register_file_0_n_105_312;
   wire execution_unit_0_register_file_0_n_105_313;
   wire execution_unit_0_register_file_0_n_105_314;
   wire execution_unit_0_register_file_0_n_105_315;
   wire execution_unit_0_register_file_0_n_105_316;
   wire execution_unit_0_register_file_0_n_105_317;
   wire execution_unit_0_register_file_0_n_105_318;
   wire execution_unit_0_register_file_0_n_105_319;
   wire execution_unit_0_register_file_0_n_106_0;
   wire execution_unit_0_register_file_0_n_106_1;
   wire execution_unit_0_register_file_0_n_106_2;
   wire execution_unit_0_register_file_0_n_106_3;
   wire execution_unit_0_register_file_0_n_106_4;
   wire execution_unit_0_register_file_0_n_106_5;
   wire execution_unit_0_register_file_0_n_106_6;
   wire execution_unit_0_register_file_0_n_106_7;
   wire execution_unit_0_register_file_0_n_106_8;
   wire execution_unit_0_register_file_0_n_106_9;
   wire execution_unit_0_register_file_0_n_106_10;
   wire execution_unit_0_register_file_0_n_106_11;
   wire execution_unit_0_register_file_0_n_106_12;
   wire execution_unit_0_register_file_0_n_106_13;
   wire [15:0]execution_unit_0_register_file_0_r1;
   wire execution_unit_0_register_file_0_n_108_0;
   wire execution_unit_0_register_file_0_n_109_0;
   wire execution_unit_0_register_file_0_n_109_1;
   wire execution_unit_0_register_file_0_n_109_2;
   wire execution_unit_0_register_file_0_n_109_3;
   wire execution_unit_0_register_file_0_n_109_4;
   wire execution_unit_0_register_file_0_n_109_5;
   wire execution_unit_0_register_file_0_n_109_6;
   wire execution_unit_0_register_file_0_n_109_7;
   wire execution_unit_0_register_file_0_n_109_8;
   wire execution_unit_0_register_file_0_n_109_9;
   wire execution_unit_0_register_file_0_n_109_10;
   wire execution_unit_0_register_file_0_n_109_11;
   wire execution_unit_0_register_file_0_n_109_12;
   wire execution_unit_0_register_file_0_n_109_13;
   wire execution_unit_0_register_file_0_n_109_14;
   wire execution_unit_0_register_file_0_n_110_0;
   wire execution_unit_0_register_file_0_n_110_1;
   wire execution_unit_0_register_file_0_n_110_2;
   wire execution_unit_0_register_file_0_n_112_0;
   wire execution_unit_0_register_file_0_n_112_1;
   wire execution_unit_0_register_file_0_n_112_2;
   wire execution_unit_0_register_file_0_n_112_3;
   wire execution_unit_0_register_file_0_n_112_4;
   wire execution_unit_0_register_file_0_n_112_5;
   wire execution_unit_0_register_file_0_n_112_6;
   wire execution_unit_0_register_file_0_n_112_7;
   wire execution_unit_0_register_file_0_n_112_8;
   wire execution_unit_0_register_file_0_n_112_9;
   wire execution_unit_0_register_file_0_n_112_10;
   wire execution_unit_0_register_file_0_n_112_11;
   wire execution_unit_0_register_file_0_n_112_12;
   wire execution_unit_0_register_file_0_n_112_13;
   wire execution_unit_0_register_file_0_n_112_14;
   wire execution_unit_0_register_file_0_n_112_15;
   wire execution_unit_0_register_file_0_n_112_16;
   wire execution_unit_0_register_file_0_n_112_17;
   wire execution_unit_0_register_file_0_n_112_18;
   wire execution_unit_0_register_file_0_n_112_19;
   wire execution_unit_0_register_file_0_n_112_20;
   wire execution_unit_0_register_file_0_n_112_21;
   wire execution_unit_0_register_file_0_n_112_22;
   wire execution_unit_0_register_file_0_n_112_23;
   wire execution_unit_0_register_file_0_n_112_24;
   wire execution_unit_0_register_file_0_n_112_25;
   wire execution_unit_0_register_file_0_n_112_26;
   wire execution_unit_0_register_file_0_n_112_27;
   wire execution_unit_0_register_file_0_n_112_28;
   wire execution_unit_0_register_file_0_n_112_29;
   wire execution_unit_0_register_file_0_n_112_30;
   wire execution_unit_0_register_file_0_n_112_31;
   wire execution_unit_0_register_file_0_n_112_32;
   wire execution_unit_0_register_file_0_n_112_33;
   wire execution_unit_0_register_file_0_n_112_34;
   wire execution_unit_0_register_file_0_n_112_35;
   wire execution_unit_0_register_file_0_n_112_36;
   wire execution_unit_0_register_file_0_n_112_37;
   wire execution_unit_0_register_file_0_n_112_38;
   wire execution_unit_0_register_file_0_n_112_39;
   wire execution_unit_0_register_file_0_n_112_40;
   wire execution_unit_0_register_file_0_n_112_41;
   wire execution_unit_0_register_file_0_n_112_42;
   wire execution_unit_0_register_file_0_n_112_43;
   wire execution_unit_0_register_file_0_n_112_44;
   wire execution_unit_0_register_file_0_n_112_45;
   wire execution_unit_0_register_file_0_n_112_46;
   wire execution_unit_0_register_file_0_n_112_47;
   wire execution_unit_0_register_file_0_n_112_48;
   wire execution_unit_0_register_file_0_n_112_49;
   wire execution_unit_0_register_file_0_n_112_50;
   wire execution_unit_0_register_file_0_n_112_51;
   wire execution_unit_0_register_file_0_n_112_52;
   wire execution_unit_0_register_file_0_n_112_53;
   wire execution_unit_0_register_file_0_n_112_54;
   wire execution_unit_0_register_file_0_n_112_55;
   wire execution_unit_0_register_file_0_n_112_56;
   wire execution_unit_0_register_file_0_n_112_57;
   wire execution_unit_0_register_file_0_n_112_58;
   wire execution_unit_0_register_file_0_n_112_59;
   wire execution_unit_0_register_file_0_n_112_60;
   wire execution_unit_0_register_file_0_n_112_61;
   wire execution_unit_0_register_file_0_n_112_62;
   wire execution_unit_0_register_file_0_n_112_63;
   wire execution_unit_0_register_file_0_n_112_64;
   wire execution_unit_0_register_file_0_n_112_65;
   wire execution_unit_0_register_file_0_n_112_66;
   wire execution_unit_0_register_file_0_n_112_67;
   wire execution_unit_0_register_file_0_n_112_68;
   wire execution_unit_0_register_file_0_n_112_69;
   wire execution_unit_0_register_file_0_n_112_70;
   wire execution_unit_0_register_file_0_n_112_71;
   wire execution_unit_0_register_file_0_n_112_72;
   wire execution_unit_0_register_file_0_n_112_73;
   wire execution_unit_0_register_file_0_n_112_74;
   wire execution_unit_0_register_file_0_n_112_75;
   wire execution_unit_0_register_file_0_n_112_76;
   wire execution_unit_0_register_file_0_n_112_77;
   wire execution_unit_0_register_file_0_n_112_78;
   wire execution_unit_0_register_file_0_n_112_79;
   wire execution_unit_0_register_file_0_n_112_80;
   wire execution_unit_0_register_file_0_n_112_81;
   wire execution_unit_0_register_file_0_n_112_82;
   wire execution_unit_0_register_file_0_n_112_83;
   wire execution_unit_0_register_file_0_n_112_84;
   wire execution_unit_0_register_file_0_n_112_85;
   wire execution_unit_0_register_file_0_n_112_86;
   wire execution_unit_0_register_file_0_n_112_87;
   wire execution_unit_0_register_file_0_n_112_88;
   wire execution_unit_0_register_file_0_n_112_89;
   wire execution_unit_0_register_file_0_n_112_90;
   wire execution_unit_0_register_file_0_n_112_91;
   wire execution_unit_0_register_file_0_n_112_92;
   wire execution_unit_0_register_file_0_n_112_93;
   wire execution_unit_0_register_file_0_n_112_94;
   wire execution_unit_0_register_file_0_n_112_95;
   wire execution_unit_0_register_file_0_n_112_96;
   wire execution_unit_0_register_file_0_n_112_97;
   wire execution_unit_0_register_file_0_n_112_98;
   wire execution_unit_0_register_file_0_n_112_99;
   wire execution_unit_0_register_file_0_n_112_100;
   wire execution_unit_0_register_file_0_n_112_101;
   wire execution_unit_0_register_file_0_n_112_102;
   wire execution_unit_0_register_file_0_n_112_103;
   wire execution_unit_0_register_file_0_n_112_104;
   wire execution_unit_0_register_file_0_n_112_105;
   wire execution_unit_0_register_file_0_n_112_106;
   wire execution_unit_0_register_file_0_n_112_107;
   wire execution_unit_0_register_file_0_n_112_108;
   wire execution_unit_0_register_file_0_n_112_109;
   wire execution_unit_0_register_file_0_n_112_110;
   wire execution_unit_0_register_file_0_n_112_111;
   wire execution_unit_0_register_file_0_n_112_112;
   wire execution_unit_0_register_file_0_n_112_113;
   wire execution_unit_0_register_file_0_n_112_114;
   wire execution_unit_0_register_file_0_n_112_115;
   wire execution_unit_0_register_file_0_n_112_116;
   wire execution_unit_0_register_file_0_n_112_117;
   wire execution_unit_0_register_file_0_n_112_118;
   wire execution_unit_0_register_file_0_n_112_119;
   wire execution_unit_0_register_file_0_n_112_120;
   wire execution_unit_0_register_file_0_n_112_121;
   wire execution_unit_0_register_file_0_n_112_122;
   wire execution_unit_0_register_file_0_n_112_123;
   wire execution_unit_0_register_file_0_n_112_124;
   wire execution_unit_0_register_file_0_n_112_125;
   wire execution_unit_0_register_file_0_n_112_126;
   wire execution_unit_0_register_file_0_n_112_127;
   wire execution_unit_0_register_file_0_n_112_128;
   wire execution_unit_0_register_file_0_n_112_129;
   wire execution_unit_0_register_file_0_n_112_130;
   wire execution_unit_0_register_file_0_n_112_131;
   wire execution_unit_0_register_file_0_n_112_132;
   wire execution_unit_0_register_file_0_n_112_133;
   wire execution_unit_0_register_file_0_n_112_134;
   wire execution_unit_0_register_file_0_n_112_135;
   wire execution_unit_0_register_file_0_n_112_136;
   wire execution_unit_0_register_file_0_n_112_137;
   wire execution_unit_0_register_file_0_n_112_138;
   wire execution_unit_0_register_file_0_n_112_139;
   wire execution_unit_0_register_file_0_n_112_140;
   wire execution_unit_0_register_file_0_n_112_141;
   wire execution_unit_0_register_file_0_n_112_142;
   wire execution_unit_0_register_file_0_n_112_143;
   wire execution_unit_0_register_file_0_n_112_144;
   wire execution_unit_0_register_file_0_n_112_145;
   wire execution_unit_0_register_file_0_n_112_146;
   wire execution_unit_0_register_file_0_n_112_147;
   wire execution_unit_0_register_file_0_n_112_148;
   wire execution_unit_0_register_file_0_n_112_149;
   wire execution_unit_0_register_file_0_n_112_150;
   wire execution_unit_0_register_file_0_n_112_151;
   wire execution_unit_0_register_file_0_n_112_152;
   wire execution_unit_0_register_file_0_n_112_153;
   wire execution_unit_0_register_file_0_n_112_154;
   wire execution_unit_0_register_file_0_n_112_155;
   wire execution_unit_0_register_file_0_n_112_156;
   wire execution_unit_0_register_file_0_n_112_157;
   wire execution_unit_0_register_file_0_n_112_158;
   wire execution_unit_0_register_file_0_n_112_159;
   wire execution_unit_0_register_file_0_n_112_160;
   wire execution_unit_0_register_file_0_n_112_161;
   wire execution_unit_0_register_file_0_n_112_162;
   wire execution_unit_0_register_file_0_n_112_163;
   wire execution_unit_0_register_file_0_n_112_164;
   wire execution_unit_0_register_file_0_n_112_165;
   wire execution_unit_0_register_file_0_n_112_166;
   wire execution_unit_0_register_file_0_n_112_167;
   wire execution_unit_0_register_file_0_n_112_168;
   wire execution_unit_0_register_file_0_n_112_169;
   wire execution_unit_0_register_file_0_n_112_170;
   wire execution_unit_0_register_file_0_n_112_171;
   wire execution_unit_0_register_file_0_n_112_172;
   wire execution_unit_0_register_file_0_n_112_173;
   wire execution_unit_0_register_file_0_n_112_174;
   wire execution_unit_0_register_file_0_n_112_175;
   wire execution_unit_0_register_file_0_n_112_176;
   wire execution_unit_0_register_file_0_n_112_177;
   wire execution_unit_0_register_file_0_n_112_178;
   wire execution_unit_0_register_file_0_n_112_179;
   wire execution_unit_0_register_file_0_n_112_180;
   wire execution_unit_0_register_file_0_n_112_181;
   wire execution_unit_0_register_file_0_n_112_182;
   wire execution_unit_0_register_file_0_n_112_183;
   wire execution_unit_0_register_file_0_n_112_184;
   wire execution_unit_0_register_file_0_n_112_185;
   wire execution_unit_0_register_file_0_n_112_186;
   wire execution_unit_0_register_file_0_n_112_187;
   wire execution_unit_0_register_file_0_n_112_188;
   wire execution_unit_0_register_file_0_n_112_189;
   wire execution_unit_0_register_file_0_n_112_190;
   wire execution_unit_0_register_file_0_n_112_191;
   wire execution_unit_0_register_file_0_n_112_192;
   wire execution_unit_0_register_file_0_n_112_193;
   wire execution_unit_0_register_file_0_n_112_194;
   wire execution_unit_0_register_file_0_n_112_195;
   wire execution_unit_0_register_file_0_n_112_196;
   wire execution_unit_0_register_file_0_n_112_197;
   wire execution_unit_0_register_file_0_n_112_198;
   wire execution_unit_0_register_file_0_n_112_199;
   wire execution_unit_0_register_file_0_n_112_200;
   wire execution_unit_0_register_file_0_n_112_201;
   wire execution_unit_0_register_file_0_n_112_202;
   wire execution_unit_0_register_file_0_n_112_203;
   wire execution_unit_0_register_file_0_n_112_204;
   wire execution_unit_0_register_file_0_n_112_205;
   wire execution_unit_0_register_file_0_n_112_206;
   wire execution_unit_0_register_file_0_n_112_207;
   wire execution_unit_0_register_file_0_n_112_208;
   wire execution_unit_0_register_file_0_n_112_209;
   wire execution_unit_0_register_file_0_n_112_210;
   wire execution_unit_0_register_file_0_n_112_211;
   wire execution_unit_0_register_file_0_n_112_212;
   wire execution_unit_0_register_file_0_n_112_213;
   wire execution_unit_0_register_file_0_n_112_214;
   wire execution_unit_0_register_file_0_n_112_215;
   wire execution_unit_0_register_file_0_n_112_216;
   wire execution_unit_0_register_file_0_n_112_217;
   wire execution_unit_0_register_file_0_n_112_218;
   wire execution_unit_0_register_file_0_n_112_219;
   wire execution_unit_0_register_file_0_n_112_220;
   wire execution_unit_0_register_file_0_n_112_221;
   wire execution_unit_0_register_file_0_n_112_222;
   wire execution_unit_0_register_file_0_n_112_223;
   wire execution_unit_0_register_file_0_n_112_224;
   wire execution_unit_0_register_file_0_n_112_225;
   wire execution_unit_0_register_file_0_n_112_226;
   wire execution_unit_0_register_file_0_n_112_227;
   wire execution_unit_0_register_file_0_n_112_228;
   wire execution_unit_0_register_file_0_n_112_229;
   wire execution_unit_0_register_file_0_n_112_230;
   wire execution_unit_0_register_file_0_n_112_231;
   wire execution_unit_0_register_file_0_n_112_232;
   wire execution_unit_0_register_file_0_n_112_233;
   wire execution_unit_0_register_file_0_n_112_234;
   wire execution_unit_0_register_file_0_n_112_235;
   wire execution_unit_0_register_file_0_n_112_236;
   wire execution_unit_0_register_file_0_n_112_237;
   wire execution_unit_0_register_file_0_n_112_238;
   wire execution_unit_0_register_file_0_n_112_239;
   wire execution_unit_0_register_file_0_n_112_240;
   wire execution_unit_0_register_file_0_n_112_241;
   wire execution_unit_0_register_file_0_n_112_242;
   wire execution_unit_0_register_file_0_n_112_243;
   wire execution_unit_0_register_file_0_n_112_244;
   wire execution_unit_0_register_file_0_n_112_245;
   wire execution_unit_0_register_file_0_n_112_246;
   wire execution_unit_0_register_file_0_n_112_247;
   wire execution_unit_0_register_file_0_n_112_248;
   wire execution_unit_0_register_file_0_n_112_249;
   wire execution_unit_0_register_file_0_n_112_250;
   wire execution_unit_0_register_file_0_n_112_251;
   wire execution_unit_0_register_file_0_n_112_252;
   wire execution_unit_0_register_file_0_n_112_253;
   wire execution_unit_0_register_file_0_n_112_254;
   wire execution_unit_0_register_file_0_n_112_255;
   wire execution_unit_0_register_file_0_n_112_256;
   wire execution_unit_0_register_file_0_n_112_257;
   wire execution_unit_0_register_file_0_n_112_258;
   wire execution_unit_0_register_file_0_n_112_259;
   wire execution_unit_0_register_file_0_n_112_260;
   wire execution_unit_0_register_file_0_n_112_261;
   wire execution_unit_0_register_file_0_n_112_262;
   wire execution_unit_0_register_file_0_n_112_263;
   wire execution_unit_0_register_file_0_n_112_264;
   wire execution_unit_0_register_file_0_n_112_265;
   wire execution_unit_0_register_file_0_n_112_266;
   wire execution_unit_0_register_file_0_n_112_267;
   wire execution_unit_0_register_file_0_n_112_268;
   wire execution_unit_0_register_file_0_n_112_269;
   wire execution_unit_0_register_file_0_n_112_270;
   wire execution_unit_0_register_file_0_n_112_271;
   wire execution_unit_0_register_file_0_n_112_272;
   wire execution_unit_0_register_file_0_n_112_273;
   wire execution_unit_0_register_file_0_n_112_274;
   wire execution_unit_0_register_file_0_n_112_275;
   wire execution_unit_0_register_file_0_n_112_276;
   wire execution_unit_0_register_file_0_n_112_277;
   wire execution_unit_0_register_file_0_n_112_278;
   wire execution_unit_0_register_file_0_n_112_279;
   wire execution_unit_0_register_file_0_n_112_280;
   wire execution_unit_0_register_file_0_n_112_281;
   wire execution_unit_0_register_file_0_n_112_282;
   wire execution_unit_0_register_file_0_n_112_283;
   wire execution_unit_0_register_file_0_n_112_284;
   wire execution_unit_0_register_file_0_n_112_285;
   wire execution_unit_0_register_file_0_n_112_286;
   wire execution_unit_0_register_file_0_n_112_287;
   wire execution_unit_0_register_file_0_n_112_288;
   wire execution_unit_0_register_file_0_n_112_289;
   wire execution_unit_0_register_file_0_n_112_290;
   wire execution_unit_0_register_file_0_n_112_291;
   wire execution_unit_0_register_file_0_n_112_292;
   wire execution_unit_0_register_file_0_n_112_293;
   wire execution_unit_0_register_file_0_n_112_294;
   wire execution_unit_0_register_file_0_n_112_295;
   wire execution_unit_0_register_file_0_n_112_296;
   wire execution_unit_0_register_file_0_n_112_297;
   wire execution_unit_0_register_file_0_n_112_298;
   wire execution_unit_0_register_file_0_n_112_299;
   wire execution_unit_0_register_file_0_n_112_300;
   wire execution_unit_0_register_file_0_n_112_301;
   wire execution_unit_0_register_file_0_n_112_302;
   wire execution_unit_0_register_file_0_n_112_303;
   wire execution_unit_0_register_file_0_n_112_304;
   wire execution_unit_0_register_file_0_n_112_305;
   wire execution_unit_0_register_file_0_n_112_306;
   wire execution_unit_0_register_file_0_n_112_307;
   wire execution_unit_0_register_file_0_n_112_308;
   wire execution_unit_0_register_file_0_n_112_309;
   wire execution_unit_0_register_file_0_n_112_310;
   wire execution_unit_0_register_file_0_n_112_311;
   wire execution_unit_0_register_file_0_n_112_312;
   wire execution_unit_0_register_file_0_n_112_313;
   wire execution_unit_0_register_file_0_n_112_314;
   wire execution_unit_0_register_file_0_n_112_315;
   wire execution_unit_0_register_file_0_n_112_316;
   wire execution_unit_0_register_file_0_n_112_317;
   wire execution_unit_0_register_file_0_n_112_318;
   wire execution_unit_0_register_file_0_n_112_319;
   wire execution_unit_0_register_file_0_n_7;
   wire execution_unit_0_register_file_0_n_17;
   wire execution_unit_0_register_file_0_n_8;
   wire execution_unit_0_register_file_0_n_16;
   wire execution_unit_0_register_file_0_n_24;
   wire execution_unit_0_register_file_0_n_22;
   wire execution_unit_0_register_file_0_n_23;
   wire execution_unit_0_register_file_0_n_21;
   wire execution_unit_0_register_file_0_n_0;
   wire execution_unit_0_register_file_0_n_272;
   wire execution_unit_0_register_file_0_n_271;
   wire execution_unit_0_register_file_0_n_41;
   wire execution_unit_0_register_file_0_n_44;
   wire execution_unit_0_register_file_0_n_27;
   wire execution_unit_0_register_file_0_n_2;
   wire execution_unit_0_register_file_0_n_39;
   wire execution_unit_0_register_file_0_n_4;
   wire execution_unit_0_register_file_0_n_37;
   wire execution_unit_0_register_file_0_n_6;
   wire execution_unit_0_register_file_0_n_35;
   wire execution_unit_0_register_file_0_n_19;
   wire execution_unit_0_register_file_0_n_33;
   wire execution_unit_0_register_file_0_n_31;
   wire execution_unit_0_register_file_0_n_25;
   wire execution_unit_0_register_file_0_n_26;
   wire execution_unit_0_register_file_0_n_29;
   wire execution_unit_0_register_file_0_n_10;
   wire execution_unit_0_register_file_0_n_14;
   wire execution_unit_0_register_file_0_n_255;
   wire execution_unit_0_register_file_0_n_273;
   wire execution_unit_0_register_file_0_n_288;
   wire execution_unit_0_register_file_0_n_270;
   wire execution_unit_0_register_file_0_n_178;
   wire execution_unit_0_register_file_0_n_181;
   wire execution_unit_0_register_file_0_n_196;
   wire execution_unit_0_register_file_0_n_179;
   wire execution_unit_0_register_file_0_n_159;
   wire execution_unit_0_register_file_0_n_162;
   wire execution_unit_0_register_file_0_n_177;
   wire execution_unit_0_register_file_0_n_160;
   wire execution_unit_0_register_file_0_n_140;
   wire execution_unit_0_register_file_0_n_143;
   wire execution_unit_0_register_file_0_n_158;
   wire execution_unit_0_register_file_0_n_141;
   wire execution_unit_0_register_file_0_n_121;
   wire execution_unit_0_register_file_0_n_124;
   wire execution_unit_0_register_file_0_n_139;
   wire execution_unit_0_register_file_0_n_122;
   wire execution_unit_0_register_file_0_n_102;
   wire execution_unit_0_register_file_0_n_105;
   wire execution_unit_0_register_file_0_n_120;
   wire execution_unit_0_register_file_0_n_103;
   wire execution_unit_0_register_file_0_n_83;
   wire execution_unit_0_register_file_0_n_86;
   wire execution_unit_0_register_file_0_n_101;
   wire execution_unit_0_register_file_0_n_84;
   wire execution_unit_0_register_file_0_n_64;
   wire execution_unit_0_register_file_0_n_67;
   wire execution_unit_0_register_file_0_n_82;
   wire execution_unit_0_register_file_0_n_65;
   wire execution_unit_0_register_file_0_n_45;
   wire execution_unit_0_register_file_0_n_48;
   wire execution_unit_0_register_file_0_n_63;
   wire execution_unit_0_register_file_0_n_46;
   wire execution_unit_0_register_file_0_n_197;
   wire execution_unit_0_register_file_0_n_200;
   wire execution_unit_0_register_file_0_n_215;
   wire execution_unit_0_register_file_0_n_198;
   wire execution_unit_0_register_file_0_n_254;
   wire execution_unit_0_register_file_0_n_235;
   wire execution_unit_0_register_file_0_n_238;
   wire execution_unit_0_register_file_0_n_253;
   wire execution_unit_0_register_file_0_n_236;
   wire execution_unit_0_register_file_0_n_216;
   wire execution_unit_0_register_file_0_n_219;
   wire execution_unit_0_register_file_0_n_234;
   wire execution_unit_0_register_file_0_n_217;
   wire execution_unit_0_register_file_0_n_28;
   wire execution_unit_0_register_file_0_n_9;
   wire execution_unit_0_register_file_0_n_13;
   wire execution_unit_0_register_file_0_n_180;
   wire execution_unit_0_register_file_0_n_161;
   wire execution_unit_0_register_file_0_n_142;
   wire execution_unit_0_register_file_0_n_123;
   wire execution_unit_0_register_file_0_n_104;
   wire execution_unit_0_register_file_0_n_85;
   wire execution_unit_0_register_file_0_n_66;
   wire execution_unit_0_register_file_0_n_47;
   wire execution_unit_0_register_file_0_n_199;
   wire execution_unit_0_register_file_0_n_237;
   wire execution_unit_0_register_file_0_n_218;
   wire execution_unit_0_register_file_0_n_30;
   wire execution_unit_0_register_file_0_n_11;
   wire execution_unit_0_register_file_0_n_15;
   wire execution_unit_0_register_file_0_n_256;
   wire execution_unit_0_register_file_0_n_274;
   wire execution_unit_0_register_file_0_n_182;
   wire execution_unit_0_register_file_0_n_163;
   wire execution_unit_0_register_file_0_n_144;
   wire execution_unit_0_register_file_0_n_125;
   wire execution_unit_0_register_file_0_n_106;
   wire execution_unit_0_register_file_0_n_87;
   wire execution_unit_0_register_file_0_n_68;
   wire execution_unit_0_register_file_0_n_49;
   wire execution_unit_0_register_file_0_n_201;
   wire execution_unit_0_register_file_0_n_239;
   wire execution_unit_0_register_file_0_n_220;
   wire execution_unit_0_register_file_0_n_257;
   wire execution_unit_0_register_file_0_n_275;
   wire execution_unit_0_register_file_0_n_183;
   wire execution_unit_0_register_file_0_n_164;
   wire execution_unit_0_register_file_0_n_145;
   wire execution_unit_0_register_file_0_n_126;
   wire execution_unit_0_register_file_0_n_107;
   wire execution_unit_0_register_file_0_n_88;
   wire execution_unit_0_register_file_0_n_69;
   wire execution_unit_0_register_file_0_n_50;
   wire execution_unit_0_register_file_0_n_202;
   wire execution_unit_0_register_file_0_n_240;
   wire execution_unit_0_register_file_0_n_221;
   wire execution_unit_0_register_file_0_n_32;
   wire execution_unit_0_register_file_0_n_258;
   wire execution_unit_0_register_file_0_n_276;
   wire execution_unit_0_register_file_0_n_184;
   wire execution_unit_0_register_file_0_n_165;
   wire execution_unit_0_register_file_0_n_146;
   wire execution_unit_0_register_file_0_n_127;
   wire execution_unit_0_register_file_0_n_108;
   wire execution_unit_0_register_file_0_n_89;
   wire execution_unit_0_register_file_0_n_70;
   wire execution_unit_0_register_file_0_n_51;
   wire execution_unit_0_register_file_0_n_203;
   wire execution_unit_0_register_file_0_n_241;
   wire execution_unit_0_register_file_0_n_222;
   wire execution_unit_0_register_file_0_n_259;
   wire execution_unit_0_register_file_0_n_277;
   wire execution_unit_0_register_file_0_n_185;
   wire execution_unit_0_register_file_0_n_166;
   wire execution_unit_0_register_file_0_n_147;
   wire execution_unit_0_register_file_0_n_128;
   wire execution_unit_0_register_file_0_n_109;
   wire execution_unit_0_register_file_0_n_90;
   wire execution_unit_0_register_file_0_n_71;
   wire execution_unit_0_register_file_0_n_52;
   wire execution_unit_0_register_file_0_n_204;
   wire execution_unit_0_register_file_0_n_242;
   wire execution_unit_0_register_file_0_n_223;
   wire execution_unit_0_register_file_0_n_34;
   wire execution_unit_0_register_file_0_n_18;
   wire execution_unit_0_register_file_0_n_260;
   wire execution_unit_0_register_file_0_n_278;
   wire execution_unit_0_register_file_0_n_186;
   wire execution_unit_0_register_file_0_n_167;
   wire execution_unit_0_register_file_0_n_148;
   wire execution_unit_0_register_file_0_n_129;
   wire execution_unit_0_register_file_0_n_110;
   wire execution_unit_0_register_file_0_n_91;
   wire execution_unit_0_register_file_0_n_72;
   wire execution_unit_0_register_file_0_n_53;
   wire execution_unit_0_register_file_0_n_205;
   wire execution_unit_0_register_file_0_n_243;
   wire execution_unit_0_register_file_0_n_224;
   wire execution_unit_0_register_file_0_n_261;
   wire execution_unit_0_register_file_0_n_279;
   wire execution_unit_0_register_file_0_n_187;
   wire execution_unit_0_register_file_0_n_168;
   wire execution_unit_0_register_file_0_n_149;
   wire execution_unit_0_register_file_0_n_130;
   wire execution_unit_0_register_file_0_n_111;
   wire execution_unit_0_register_file_0_n_92;
   wire execution_unit_0_register_file_0_n_73;
   wire execution_unit_0_register_file_0_n_54;
   wire execution_unit_0_register_file_0_n_206;
   wire execution_unit_0_register_file_0_n_244;
   wire execution_unit_0_register_file_0_n_225;
   wire execution_unit_0_register_file_0_n_36;
   wire execution_unit_0_register_file_0_n_12;
   wire execution_unit_0_register_file_0_n_20;
   wire execution_unit_0_register_file_0_n_262;
   wire execution_unit_0_register_file_0_n_280;
   wire execution_unit_0_register_file_0_n_188;
   wire execution_unit_0_register_file_0_n_169;
   wire execution_unit_0_register_file_0_n_150;
   wire execution_unit_0_register_file_0_n_131;
   wire execution_unit_0_register_file_0_n_112;
   wire execution_unit_0_register_file_0_n_93;
   wire execution_unit_0_register_file_0_n_74;
   wire execution_unit_0_register_file_0_n_55;
   wire execution_unit_0_register_file_0_n_207;
   wire execution_unit_0_register_file_0_n_245;
   wire execution_unit_0_register_file_0_n_226;
   wire execution_unit_0_register_file_0_n_263;
   wire execution_unit_0_register_file_0_n_281;
   wire execution_unit_0_register_file_0_n_189;
   wire execution_unit_0_register_file_0_n_170;
   wire execution_unit_0_register_file_0_n_151;
   wire execution_unit_0_register_file_0_n_132;
   wire execution_unit_0_register_file_0_n_113;
   wire execution_unit_0_register_file_0_n_94;
   wire execution_unit_0_register_file_0_n_75;
   wire execution_unit_0_register_file_0_n_56;
   wire execution_unit_0_register_file_0_n_208;
   wire execution_unit_0_register_file_0_n_246;
   wire execution_unit_0_register_file_0_n_227;
   wire execution_unit_0_register_file_0_n_38;
   wire execution_unit_0_register_file_0_n_5;
   wire execution_unit_0_register_file_0_n_264;
   wire execution_unit_0_register_file_0_n_282;
   wire execution_unit_0_register_file_0_n_190;
   wire execution_unit_0_register_file_0_n_171;
   wire execution_unit_0_register_file_0_n_152;
   wire execution_unit_0_register_file_0_n_133;
   wire execution_unit_0_register_file_0_n_114;
   wire execution_unit_0_register_file_0_n_95;
   wire execution_unit_0_register_file_0_n_76;
   wire execution_unit_0_register_file_0_n_57;
   wire execution_unit_0_register_file_0_n_209;
   wire execution_unit_0_register_file_0_n_247;
   wire execution_unit_0_register_file_0_n_228;
   wire execution_unit_0_register_file_0_n_265;
   wire execution_unit_0_register_file_0_n_283;
   wire execution_unit_0_register_file_0_n_191;
   wire execution_unit_0_register_file_0_n_172;
   wire execution_unit_0_register_file_0_n_153;
   wire execution_unit_0_register_file_0_n_134;
   wire execution_unit_0_register_file_0_n_115;
   wire execution_unit_0_register_file_0_n_96;
   wire execution_unit_0_register_file_0_n_77;
   wire execution_unit_0_register_file_0_n_58;
   wire execution_unit_0_register_file_0_n_210;
   wire execution_unit_0_register_file_0_n_248;
   wire execution_unit_0_register_file_0_n_229;
   wire execution_unit_0_register_file_0_n_40;
   wire execution_unit_0_register_file_0_n_3;
   wire execution_unit_0_register_file_0_n_266;
   wire execution_unit_0_register_file_0_n_284;
   wire execution_unit_0_register_file_0_n_192;
   wire execution_unit_0_register_file_0_n_173;
   wire execution_unit_0_register_file_0_n_154;
   wire execution_unit_0_register_file_0_n_135;
   wire execution_unit_0_register_file_0_n_116;
   wire execution_unit_0_register_file_0_n_97;
   wire execution_unit_0_register_file_0_n_78;
   wire execution_unit_0_register_file_0_n_59;
   wire execution_unit_0_register_file_0_n_211;
   wire execution_unit_0_register_file_0_n_249;
   wire execution_unit_0_register_file_0_n_230;
   wire execution_unit_0_register_file_0_n_267;
   wire execution_unit_0_register_file_0_n_285;
   wire execution_unit_0_register_file_0_n_193;
   wire execution_unit_0_register_file_0_n_174;
   wire execution_unit_0_register_file_0_n_155;
   wire execution_unit_0_register_file_0_n_136;
   wire execution_unit_0_register_file_0_n_117;
   wire execution_unit_0_register_file_0_n_98;
   wire execution_unit_0_register_file_0_n_79;
   wire execution_unit_0_register_file_0_n_60;
   wire execution_unit_0_register_file_0_n_212;
   wire execution_unit_0_register_file_0_n_250;
   wire execution_unit_0_register_file_0_n_231;
   wire execution_unit_0_register_file_0_n_42;
   wire execution_unit_0_register_file_0_n_1;
   wire execution_unit_0_register_file_0_n_268;
   wire execution_unit_0_register_file_0_n_286;
   wire execution_unit_0_register_file_0_n_194;
   wire execution_unit_0_register_file_0_n_175;
   wire execution_unit_0_register_file_0_n_156;
   wire execution_unit_0_register_file_0_n_137;
   wire execution_unit_0_register_file_0_n_118;
   wire execution_unit_0_register_file_0_n_99;
   wire execution_unit_0_register_file_0_n_80;
   wire execution_unit_0_register_file_0_n_61;
   wire execution_unit_0_register_file_0_n_213;
   wire execution_unit_0_register_file_0_n_251;
   wire execution_unit_0_register_file_0_n_232;
   wire execution_unit_0_register_file_0_n_269;
   wire execution_unit_0_register_file_0_n_287;
   wire execution_unit_0_register_file_0_n_195;
   wire execution_unit_0_register_file_0_n_176;
   wire execution_unit_0_register_file_0_n_157;
   wire execution_unit_0_register_file_0_n_138;
   wire execution_unit_0_register_file_0_n_119;
   wire execution_unit_0_register_file_0_n_100;
   wire execution_unit_0_register_file_0_n_81;
   wire execution_unit_0_register_file_0_n_62;
   wire execution_unit_0_register_file_0_n_214;
   wire execution_unit_0_register_file_0_n_252;
   wire execution_unit_0_register_file_0_n_233;
   wire execution_unit_0_register_file_0_n_43;
   wire clock_module_0_cpuoff_and_mclk_dma_wkup;
   wire clock_module_0_cpuoff_and_mclk_dma_wkup_s;
   wire clock_module_0_mclk_wkup_s;
   wire clock_module_0_cpuoff_and_mclk_dma_enable;
   wire clock_module_0_por_noscan;
   wire clock_module_0_puc_a_scan;
   wire clock_module_0_puc_noscan_n;
   wire clock_module_0_scg0_and_mclk_dma_enable;
   wire clock_module_0_cpuoff_and_mclk_enable;
   wire clock_module_0_cpu_enabled_with_dco;
   wire clock_module_0_dco_not_enabled_by_dbg;
   wire clock_module_0_dco_disable_by_scg0;
   wire clock_module_0_dco_disable_by_cpu_en;
   wire clock_module_0_dco_enable_nxt;
   wire clock_module_0_scg0_and_mclk_dma_wkup;
   wire clock_module_0_dco_en_wkup;
   wire clock_module_0_dco_mclk_wkup;
   wire clock_module_0_dco_wkup_set_scan_observe;
   wire clock_module_0_dco_wkup_set_scan;
   wire clock_module_0_dco_wkup_n;
   wire clock_module_0_scg1_and_mclk_dma_enable;
   wire clock_module_0_scg1_and_mclk_dma_wkup;
   wire clock_module_0_scg1_and_mclk_dma_wkup_s;
   wire clock_module_0_nodiv_mclk_n;
   wire clock_module_0_dco_disable;
   wire clock_module_0_n_1_0;
   wire clock_module_0_n_7_0;
   wire clock_module_0_n_7_1;
   wire clock_module_0_n_7_2;
   wire clock_module_0_n_7_3;
   wire clock_module_0_reg_sel;
   wire clock_module_0_reg_read;
   wire clock_module_0_n_10_0;
   wire clock_module_0_n_11_0;
   wire clock_module_0_reg_lo_write;
   wire clock_module_0_bcsctl2_wr;
   wire [7:0]clock_module_0_bcsctl2;
   wire clock_module_0_reg_hi_write;
   wire clock_module_0_bcsctl1_wr;
   wire [7:0]clock_module_0_bcsctl1;
   wire [2:0]clock_module_0_aclk_div;
   wire clock_module_0_n_23_0;
   wire clock_module_0_n_23_1;
   wire clock_module_0_n_28_0;
   wire clock_module_0_n_28_1;
   wire clock_module_0_n_28_2;
   wire clock_module_0_n_28_3;
   wire clock_module_0_n_28_4;
   wire clock_module_0_n_28_5;
   wire clock_module_0_n_28_6;
   wire clock_module_0_n_28_7;
   wire clock_module_0_n_28_8;
   wire clock_module_0_n_28_9;
   wire clock_module_0_aclk_div_sel;
   wire clock_module_0_n_29_0;
   wire clock_module_0_aclk_div_en;
   wire [2:0]clock_module_0_mclk_div;
   wire clock_module_0_n_31_0;
   wire clock_module_0_n_31_1;
   wire clock_module_0_n_36_0;
   wire clock_module_0_n_36_1;
   wire clock_module_0_n_36_2;
   wire clock_module_0_n_36_3;
   wire clock_module_0_n_36_4;
   wire clock_module_0_n_36_5;
   wire clock_module_0_n_36_6;
   wire clock_module_0_n_36_7;
   wire clock_module_0_n_36_8;
   wire clock_module_0_n_36_9;
   wire clock_module_0_mclk_div_sel;
   wire clock_module_0_n_37_0;
   wire clock_module_0_n_37_1;
   wire clock_module_0_mclk_active;
   wire clock_module_0_mclk_div_en;
   wire clock_module_0_n_39_0;
   wire clock_module_0_mclk_dma_div_en;
   wire clock_module_0_por_a;
   wire clock_module_0_dbg_rst_nxt;
   wire clock_module_0_dbg_rst_noscan;
   wire clock_module_0_dco_wkup_set;
   wire clock_module_0_n_46_0;
   wire [2:0]clock_module_0_smclk_div;
   wire clock_module_0_n_48_0;
   wire clock_module_0_n_48_1;
   wire clock_module_0_n_53_0;
   wire clock_module_0_n_53_1;
   wire clock_module_0_n_53_2;
   wire clock_module_0_n_53_3;
   wire clock_module_0_n_53_4;
   wire clock_module_0_n_53_5;
   wire clock_module_0_n_53_6;
   wire clock_module_0_n_53_7;
   wire clock_module_0_n_53_8;
   wire clock_module_0_n_53_9;
   wire clock_module_0_smclk_div_sel;
   wire clock_module_0_n_54_0;
   wire clock_module_0_n_54_1;
   wire clock_module_0_n_54_2;
   wire clock_module_0_smclk_div_en;
   wire clock_module_0_puc_a;
   wire clock_module_0_n_5;
   wire clock_module_0_n_4;
   wire clock_module_0_n_8;
   wire clock_module_0_n_10;
   wire clock_module_0_n_19;
   wire clock_module_0_n_22;
   wire clock_module_0_n_18;
   wire clock_module_0_n_20;
   wire clock_module_0_n_21;
   wire clock_module_0_n_23;
   wire clock_module_0_n_24;
   wire clock_module_0_n_1;
   wire clock_module_0_n_28;
   wire clock_module_0_n_9;
   wire clock_module_0_n_12;
   wire clock_module_0_n_15;
   wire clock_module_0_n_11;
   wire clock_module_0_n_13;
   wire clock_module_0_n_14;
   wire clock_module_0_n_16;
   wire clock_module_0_n_17;
   wire clock_module_0_n_39;
   wire clock_module_0_n_38;
   wire clock_module_0_n_40;
   wire clock_module_0_n_25;
   wire clock_module_0_n_36;
   wire clock_module_0_n_37;
   wire clock_module_0_n_26;
   wire clock_module_0_n_0;
   wire clock_module_0_n_2;
   wire clock_module_0_n_41;
   wire clock_module_0_n_27;
   wire clock_module_0_n_3;
   wire clock_module_0_n_6;
   wire clock_module_0_n_7;
   wire clock_module_0_n_30;
   wire clock_module_0_n_33;
   wire clock_module_0_n_29;
   wire clock_module_0_n_31;
   wire clock_module_0_n_32;
   wire clock_module_0_n_34;
   wire clock_module_0_n_35;
   wire clock_module_0_sync_cell_mclk_wkup_n_0;
   wire clock_module_0_sync_cell_mclk_wkup_n_1;
   wire clock_module_0_clock_gate_mclk_enable_in;
   wire clock_module_0_clock_gate_mclk_enable_latch;
   wire clock_module_0_clock_gate_mclk_n_0;
   wire clock_module_0_sync_reset_por_n_0;
   wire clock_module_0_sync_reset_por_n_1;
   wire clock_module_0_scan_mux_por_n_0_0;
   wire clock_module_0_scan_mux_por_n_0_1;
   wire clock_module_0_scan_mux_puc_rst_a_n_0_0;
   wire clock_module_0_scan_mux_puc_rst_a_n_0_1;
   wire clock_module_0_sync_cell_puc_n_0;
   wire clock_module_0_sync_cell_puc_n_1;
   wire clock_module_0_scan_mux_puc_rst_n_0_0;
   wire clock_module_0_scan_mux_puc_rst_n_0_1;
   wire clock_module_0_sync_cell_mclk_dma_wkup_n_0;
   wire clock_module_0_sync_cell_mclk_dma_wkup_n_1;
   wire clock_module_0_clock_gate_dma_mclk_enable_in;
   wire clock_module_0_clock_gate_dma_mclk_enable_latch;
   wire clock_module_0_clock_gate_dma_mclk_n_0;
   wire clock_module_0_clock_gate_aclk_enable_in;
   wire clock_module_0_clock_gate_aclk_enable_latch;
   wire clock_module_0_clock_gate_aclk_n_0;
   wire clock_module_0_clock_gate_dbg_clk_enable_in;
   wire clock_module_0_clock_gate_dbg_clk_enable_latch;
   wire clock_module_0_clock_gate_dbg_clk_n_0;
   wire clock_module_0_scan_mux_dbg_rst_n_0_0;
   wire clock_module_0_scan_mux_dbg_rst_n_0_1;
   wire clock_module_0_scan_mux_dco_wkup_observe_n_0_0;
   wire clock_module_0_scan_mux_dco_wkup_observe_n_0_1;
   wire clock_module_0_scan_mux_dco_wkup_n_0_0;
   wire clock_module_0_scan_mux_dco_wkup_n_0_1;
   wire clock_module_0_sync_cell_dco_wkup_n_0;
   wire clock_module_0_sync_cell_dco_wkup_n_1;
   wire clock_module_0_sync_cell_smclk_dma_wkup_n_0;
   wire clock_module_0_sync_cell_smclk_dma_wkup_n_1;
   wire clock_module_0_clock_gate_smclk_enable_in;
   wire clock_module_0_clock_gate_smclk_enable_latch;
   wire clock_module_0_clock_gate_smclk_n_0;
  assign per_dout_wdog[15] = 1'b0;
  assign per_dout_wdog[14] = per_dout_wdog[5];
  assign per_dout_wdog[13] = per_dout_wdog[5];
  assign per_dout_wdog[12] = 1'b0;
  assign per_dout_wdog[11] = per_dout_wdog[5];
  assign per_dout_wdog[10] = 1'b0;
  assign per_dout_wdog[9] = 1'b0;
  assign per_dout_wdog[8] = per_dout_wdog[5];
  assign cpu_id[31] = 1'b0;
  assign cpu_id[30] = 1'b0;
  assign cpu_id[29] = 1'b0;
  assign cpu_id[28] = 1'b1;
  assign cpu_id[27] = 1'b0;
  assign cpu_id[26] = 1'b0;
  assign cpu_id[25] = 1'b0;
  assign cpu_id[24] = 1'b0;
  assign cpu_id[23] = 1'b0;
  assign cpu_id[22] = 1'b0;
  assign cpu_id[21] = 1'b0;
  assign cpu_id[20] = 1'b1;
  assign cpu_id[19] = 1'b0;
  assign cpu_id[18] = 1'b0;
  assign cpu_id[17] = 1'b0;
  assign cpu_id[16] = 1'b1;
  assign cpu_id[15] = 1'b0;
  assign cpu_id[14] = 1'b0;
  assign cpu_id[13] = 1'b0;
  assign cpu_id[12] = 1'b0;
  assign cpu_id[11] = 1'b0;
  assign cpu_id[10] = 1'b0;
  assign cpu_id[9] = 1'b1;
  assign cpu_id[8] = 1'b0;
  assign cpu_id[7] = 1'b0;
  assign cpu_id[6] = 1'b0;
  assign cpu_id[5] = 1'b0;
  assign cpu_id[4] = 1'b0;
  assign cpu_id[3] = 1'b1;
  assign cpu_id[2] = 1'b0;
  assign cpu_id[1] = 1'b1;
  assign cpu_id[0] = 1'b1;
  assign dbg_i2c_sda_out = 1'b1;
  assign per_addr[13] = 1'b0;
  assign per_addr[12] = 1'b0;
  assign per_addr[11] = 1'b0;
  assign per_addr[10] = 1'b0;
  assign per_addr[9] = 1'b0;
  assign per_addr[8] = 1'b0;
  assign n_14 = pc_nxt[15];
  assign n_13 = pc_nxt[14];
  assign n_12 = pc_nxt[13];
  assign n_11 = pc_nxt[12];
  assign n_10 = pc_nxt[11];
  assign n_9 = pc_nxt[10];
  assign n_8 = pc_nxt[9];
  assign n_7 = pc_nxt[8];
  assign n_6 = pc_nxt[7];
  assign n_5 = pc_nxt[6];
  assign n_4 = pc_nxt[5];
  assign n_3 = pc_nxt[4];
  assign n_2 = pc_nxt[3];
  assign n_1 = pc_nxt[2];
  assign n_0 = pc_nxt[1];
  assign uc_0 = pc_nxt[0];
  assign execution_unit_0_alu_stat_wr[3] = execution_unit_0_alu_stat_wr[0];
  assign execution_unit_0_alu_stat_wr[2] = execution_unit_0_alu_stat_wr[0];
  assign execution_unit_0_alu_stat_wr[1] = execution_unit_0_alu_stat_wr[0];
  assign pc_sw[7] = execution_unit_0_alu_out[7];
  assign pc_sw[6] = execution_unit_0_alu_out[6];
  assign pc_sw[5] = execution_unit_0_alu_out[5];
  assign pc_sw[4] = execution_unit_0_alu_out[4];
  assign pc_sw[3] = execution_unit_0_alu_out[3];
  assign pc_sw[2] = execution_unit_0_alu_out[2];
  assign pc_sw[1] = execution_unit_0_alu_out[1];
  assign pc_sw[0] = execution_unit_0_alu_out[0];
  assign cpu_en_s = cpu_en;
  assign dbg_en_s = dbg_en;
  assign aclk_en = 1'b1;
  assign lfxt_enable = 1'b1;
  assign lfxt_wkup = 1'b0;
  assign smclk_en = 1'b1;
  NOR2_X1_LVT watchdog_0_i_1_0 (.ZN(watchdog_0_n_1), .A1(per_we[0]), .A2(
      per_we[1]));
  NAND3_X1_LVT watchdog_0_i_0_0 (.ZN(watchdog_0_n_0_0), .A1(per_addr[4]), .A2(
      per_addr[7]), .A3(per_en));
  NOR4_X1_LVT watchdog_0_i_0_1 (.ZN(watchdog_0_n_0_1), .A1(watchdog_0_n_0_0), 
      .A2(per_addr[12]), .A3(per_addr[13]), .A4(per_addr[0]));
  NOR4_X1_LVT watchdog_0_i_0_2 (.ZN(watchdog_0_n_0_2), .A1(per_addr[2]), .A2(
      per_addr[3]), .A3(per_addr[5]), .A4(per_addr[6]));
  NOR4_X1_LVT watchdog_0_i_0_3 (.ZN(watchdog_0_n_0_3), .A1(per_addr[8]), .A2(
      per_addr[9]), .A3(per_addr[10]), .A4(per_addr[11]));
  NAND3_X1_LVT watchdog_0_i_0_4 (.ZN(watchdog_0_n_0_4), .A1(watchdog_0_n_0_1), 
      .A2(watchdog_0_n_0_2), .A3(watchdog_0_n_0_3));
  NOR2_X1_LVT watchdog_0_i_0_5 (.ZN(watchdog_0_n_0), .A1(watchdog_0_n_0_4), .A2(
      per_addr[1]));
  AND2_X1_LVT watchdog_0_i_2_0 (.ZN(per_dout_wdog[5]), .A1(watchdog_0_n_1), .A2(
      watchdog_0_n_0));
  OR2_X1_LVT watchdog_0_i_3_0 (.ZN(watchdog_0_n_2), .A1(per_we[0]), .A2(per_we[1]));
  AND2_X1_LVT watchdog_0_i_4_0 (.ZN(watchdog_0_reg_wr), .A1(watchdog_0_n_2), .A2(
      watchdog_0_n_0));
  CLKGATETST_X1_LVT watchdog_0_clk_gate_wdtctl_reg (.GCK(watchdog_0_n_3), .CK(
      mclk), .E(watchdog_0_reg_wr), .SE(1'b0));
  INV_X1_LVT watchdog_0_i_5_0 (.ZN(watchdog_0_n_4), .A(puc_rst));
  DFFR_X1_LVT \watchdog_0_wdtctl_reg[7] (.Q(watchdog_0_wdtctl[7]), .QN(), .CK(
      watchdog_0_n_3), .D(per_din[7]), .RN(watchdog_0_n_4));
  AND2_X1_LVT watchdog_0_i_7_6 (.ZN(per_dout_wdog[7]), .A1(per_dout_wdog[5]), 
      .A2(watchdog_0_wdtctl[7]));
  DFFR_X1_LVT \watchdog_0_wdtctl_reg[6] (.Q(wdtnmies), .QN(), .CK(watchdog_0_n_3), 
      .D(per_din[6]), .RN(watchdog_0_n_4));
  AND2_X1_LVT watchdog_0_i_7_5 (.ZN(per_dout_wdog[6]), .A1(per_dout_wdog[5]), 
      .A2(wdtnmies));
  DFFR_X1_LVT \watchdog_0_wdtctl_reg[4] (.Q(watchdog_0_wdtctl[4]), .QN(), .CK(
      watchdog_0_n_3), .D(per_din[4]), .RN(watchdog_0_n_4));
  AND2_X1_LVT watchdog_0_i_7_4 (.ZN(per_dout_wdog[4]), .A1(per_dout_wdog[5]), 
      .A2(watchdog_0_wdtctl[4]));
  DFFR_X1_LVT \watchdog_0_wdtctl_reg[3] (.Q(watchdog_0_wdtctl[3]), .QN(), .CK(
      watchdog_0_n_3), .D(1'b0), .RN(watchdog_0_n_4));
  AND2_X1_LVT watchdog_0_i_7_3 (.ZN(per_dout_wdog[3]), .A1(per_dout_wdog[5]), 
      .A2(watchdog_0_wdtctl[3]));
  DFFR_X1_LVT \watchdog_0_wdtctl_reg[2] (.Q(watchdog_0_wdtctl[2]), .QN(), .CK(
      watchdog_0_n_3), .D(1'b0), .RN(watchdog_0_n_4));
  AND2_X1_LVT watchdog_0_i_7_2 (.ZN(per_dout_wdog[2]), .A1(per_dout_wdog[5]), 
      .A2(watchdog_0_wdtctl[2]));
  DFFR_X1_LVT \watchdog_0_wdtctl_reg[1] (.Q(watchdog_0_wdtctl[1]), .QN(), .CK(
      watchdog_0_n_3), .D(per_din[1]), .RN(watchdog_0_n_4));
  AND2_X1_LVT watchdog_0_i_7_1 (.ZN(per_dout_wdog[1]), .A1(per_dout_wdog[5]), 
      .A2(watchdog_0_wdtctl[1]));
  DFFR_X1_LVT \watchdog_0_wdtctl_reg[0] (.Q(watchdog_0_wdtctl[0]), .QN(), .CK(
      watchdog_0_n_3), .D(per_din[0]), .RN(watchdog_0_n_4));
  AND2_X1_LVT watchdog_0_i_7_0 (.ZN(per_dout_wdog[0]), .A1(watchdog_0_wdtctl[0]), 
      .A2(per_dout_wdog[5]));
  INV_X1_LVT watchdog_0_i_32_0 (.ZN(watchdog_0_n_30), .A(
      watchdog_0_wdt_evt_toggle));
  INV_X1_LVT watchdog_0_sync_reset_por_i_0_0 (.ZN(watchdog_0_sync_reset_por_n_0), 
      .A(puc_rst));
  DFFS_X1_LVT \watchdog_0_sync_reset_por_data_sync_reg[0] (.Q(
      watchdog_0_sync_reset_por_n_1), .QN(), .CK(smclk), .D(1'b0), .SN(
      watchdog_0_sync_reset_por_n_0));
  DFFS_X1_LVT \watchdog_0_sync_reset_por_data_sync_reg[1] (.Q(
      watchdog_0_wdt_rst_noscan), .QN(), .CK(smclk), .D(
      watchdog_0_sync_reset_por_n_1), .SN(watchdog_0_sync_reset_por_n_0));
  INV_X1_LVT watchdog_0_scan_mux_wdt_rst_i_0_0 (.ZN(
      watchdog_0_scan_mux_wdt_rst_n_0_0), .A(scan_mode));
  AOI22_X1_LVT watchdog_0_scan_mux_wdt_rst_i_0_1 (.ZN(
      watchdog_0_scan_mux_wdt_rst_n_0_1), .A1(watchdog_0_scan_mux_wdt_rst_n_0_0), 
      .A2(watchdog_0_wdt_rst_noscan), .B1(puc_rst), .B2(scan_mode));
  INV_X1_LVT watchdog_0_scan_mux_wdt_rst_i_0_2 (.ZN(watchdog_0_wdt_rst), .A(
      watchdog_0_scan_mux_wdt_rst_n_0_1));
  INV_X1_LVT watchdog_0_i_30_0 (.ZN(watchdog_0_n_29), .A(watchdog_0_wdt_rst));
  DFFR_X1_LVT \watchdog_0_wdtisx_s_reg[0] (.Q(watchdog_0_wdtisx_s[0]), .QN(), .CK(
      smclk), .D(watchdog_0_wdtctl[0]), .RN(watchdog_0_n_29));
  DFFR_X1_LVT \watchdog_0_wdtisx_ss_reg[0] (.Q(watchdog_0_wdtisx_ss[0]), .QN(), 
      .CK(smclk), .D(watchdog_0_wdtisx_s[0]), .RN(watchdog_0_n_29));
  INV_X1_LVT watchdog_0_i_28_0 (.ZN(watchdog_0_n_28_0), .A(
      watchdog_0_wdtisx_ss[0]));
  DFFR_X1_LVT \watchdog_0_wdtisx_s_reg[1] (.Q(watchdog_0_wdtisx_s[1]), .QN(), 
      .CK(smclk), .D(watchdog_0_wdtctl[1]), .RN(watchdog_0_n_29));
  DFFR_X1_LVT \watchdog_0_wdtisx_ss_reg[1] (.Q(watchdog_0_wdtisx_ss[1]), .QN(), 
      .CK(smclk), .D(watchdog_0_wdtisx_s[1]), .RN(watchdog_0_n_29));
  AND2_X1_LVT watchdog_0_i_28_1 (.ZN(watchdog_0_n_28_1), .A1(watchdog_0_n_28_0), 
      .A2(watchdog_0_wdtisx_ss[1]));
  NOR2_X1_LVT watchdog_0_i_28_2 (.ZN(watchdog_0_n_28_2), .A1(watchdog_0_n_28_0), 
      .A2(watchdog_0_wdtisx_ss[1]));
  NOR2_X1_LVT watchdog_0_i_28_3 (.ZN(watchdog_0_n_28_3), .A1(
      watchdog_0_wdtisx_ss[0]), .A2(watchdog_0_wdtisx_ss[1]));
  INV_X1_LVT watchdog_0_i_40_0 (.ZN(watchdog_0_n_35), .A(
      watchdog_0_wdtcnt_clr_toggle));
  AND2_X1_LVT watchdog_0_i_38_0 (.ZN(watchdog_0_wdtcnt_clr_detect), .A1(
      per_din[3]), .A2(watchdog_0_reg_wr));
  CLKGATETST_X1_LVT watchdog_0_clk_gate_wdtcnt_clr_toggle_reg (.GCK(
      watchdog_0_n_34), .CK(mclk), .E(watchdog_0_wdtcnt_clr_detect), .SE(1'b0));
  DFFR_X1_LVT watchdog_0_wdtcnt_clr_toggle_reg (.Q(watchdog_0_wdtcnt_clr_toggle), 
      .QN(), .CK(watchdog_0_n_34), .D(watchdog_0_n_35), .RN(watchdog_0_n_4));
  INV_X1_LVT watchdog_0_sync_cell_wdtcnt_clr_i_0_0 (.ZN(
      watchdog_0_sync_cell_wdtcnt_clr_n_0), .A(watchdog_0_wdt_rst));
  DFFR_X1_LVT \watchdog_0_sync_cell_wdtcnt_clr_data_sync_reg[0] (.Q(
      watchdog_0_sync_cell_wdtcnt_clr_n_1), .QN(), .CK(smclk), .D(
      watchdog_0_wdtcnt_clr_toggle), .RN(watchdog_0_sync_cell_wdtcnt_clr_n_0));
  DFFR_X1_LVT \watchdog_0_sync_cell_wdtcnt_clr_data_sync_reg[1] (.Q(
      watchdog_0_wdtcnt_clr_sync), .QN(), .CK(smclk), .D(
      watchdog_0_sync_cell_wdtcnt_clr_n_1), .RN(
      watchdog_0_sync_cell_wdtcnt_clr_n_0));
  DFFR_X1_LVT watchdog_0_wdtcnt_clr_sync_dly_reg (.Q(
      watchdog_0_wdtcnt_clr_sync_dly), .QN(), .CK(smclk), .D(
      watchdog_0_wdtcnt_clr_sync), .RN(watchdog_0_n_29));
  XOR2_X1_LVT watchdog_0_i_19_0 (.Z(watchdog_0_n_19_0), .A(
      watchdog_0_wdtcnt_clr_sync), .B(watchdog_0_wdtcnt_clr_sync_dly));
  OR2_X1_LVT watchdog_0_i_19_1 (.ZN(watchdog_0_wdtcnt_clr), .A1(
      watchdog_0_n_19_0), .A2(watchdog_0_wdtqn_edge));
  INV_X1_LVT watchdog_0_i_21_0 (.ZN(watchdog_0_n_21_0), .A(watchdog_0_wdtcnt_clr));
  AND2_X1_LVT watchdog_0_i_21_7 (.ZN(watchdog_0_n_17), .A1(watchdog_0_n_21_0), 
      .A2(watchdog_0_wdtcnt_nxt[6]));
  INV_X1_LVT watchdog_0_i_34_0 (.ZN(watchdog_0_n_31), .A(watchdog_0_wdtctl[7]));
  INV_X1_LVT watchdog_0_i_37_0 (.ZN(watchdog_0_n_37_0), .A(watchdog_0_n_31));
  NOR2_X1_LVT watchdog_0_i_37_1 (.ZN(watchdog_0_n_33), .A1(watchdog_0_n_37_0), 
      .A2(dbg_freeze));
  INV_X1_LVT watchdog_0_sync_cell_wdtcnt_incr_i_0_0 (.ZN(
      watchdog_0_sync_cell_wdtcnt_incr_n_0), .A(watchdog_0_wdt_rst));
  DFFR_X1_LVT \watchdog_0_sync_cell_wdtcnt_incr_data_sync_reg[0] (.Q(
      watchdog_0_sync_cell_wdtcnt_incr_n_1), .QN(), .CK(smclk), .D(
      watchdog_0_n_33), .RN(watchdog_0_sync_cell_wdtcnt_incr_n_0));
  DFFR_X1_LVT \watchdog_0_sync_cell_wdtcnt_incr_data_sync_reg[1] (.Q(
      watchdog_0_wdtcnt_incr), .QN(), .CK(smclk), .D(
      watchdog_0_sync_cell_wdtcnt_incr_n_1), .RN(
      watchdog_0_sync_cell_wdtcnt_incr_n_0));
  INV_X1_LVT watchdog_0_i_22_1 (.ZN(watchdog_0_n_22_1), .A(
      watchdog_0_wdtcnt_incr));
  INV_X1_LVT watchdog_0_i_22_0 (.ZN(watchdog_0_n_22_0), .A(watchdog_0_wdtcnt_clr));
  NAND2_X1_LVT watchdog_0_i_22_2 (.ZN(watchdog_0_n_27), .A1(watchdog_0_n_22_1), 
      .A2(watchdog_0_n_22_0));
  CLKGATETST_X1_LVT watchdog_0_clk_gate_wdtcnt_reg (.GCK(watchdog_0_n_10), .CK(
      smclk), .E(watchdog_0_n_27), .SE(1'b0));
  DFFR_X1_LVT \watchdog_0_wdtcnt_reg[6] (.Q(watchdog_0_wdtcnt[6]), .QN(), .CK(
      watchdog_0_n_10), .D(watchdog_0_n_17), .RN(watchdog_0_n_29));
  AND2_X1_LVT watchdog_0_i_21_6 (.ZN(watchdog_0_n_16), .A1(watchdog_0_n_21_0), 
      .A2(watchdog_0_wdtcnt_nxt[5]));
  DFFR_X1_LVT \watchdog_0_wdtcnt_reg[5] (.Q(watchdog_0_wdtcnt[5]), .QN(), .CK(
      watchdog_0_n_10), .D(watchdog_0_n_16), .RN(watchdog_0_n_29));
  AND2_X1_LVT watchdog_0_i_21_5 (.ZN(watchdog_0_n_15), .A1(watchdog_0_n_21_0), 
      .A2(watchdog_0_wdtcnt_nxt[4]));
  DFFR_X1_LVT \watchdog_0_wdtcnt_reg[4] (.Q(watchdog_0_wdtcnt[4]), .QN(), .CK(
      watchdog_0_n_10), .D(watchdog_0_n_15), .RN(watchdog_0_n_29));
  AND2_X1_LVT watchdog_0_i_21_4 (.ZN(watchdog_0_n_14), .A1(watchdog_0_n_21_0), 
      .A2(watchdog_0_wdtcnt_nxt[3]));
  DFFR_X1_LVT \watchdog_0_wdtcnt_reg[3] (.Q(watchdog_0_wdtcnt[3]), .QN(), .CK(
      watchdog_0_n_10), .D(watchdog_0_n_14), .RN(watchdog_0_n_29));
  AND2_X1_LVT watchdog_0_i_21_3 (.ZN(watchdog_0_n_13), .A1(watchdog_0_n_21_0), 
      .A2(watchdog_0_wdtcnt_nxt[2]));
  DFFR_X1_LVT \watchdog_0_wdtcnt_reg[2] (.Q(watchdog_0_wdtcnt[2]), .QN(), .CK(
      watchdog_0_n_10), .D(watchdog_0_n_13), .RN(watchdog_0_n_29));
  AND2_X1_LVT watchdog_0_i_21_2 (.ZN(watchdog_0_n_12), .A1(watchdog_0_n_21_0), 
      .A2(watchdog_0_wdtcnt_nxt[1]));
  DFFR_X1_LVT \watchdog_0_wdtcnt_reg[1] (.Q(watchdog_0_wdtcnt[1]), .QN(), .CK(
      watchdog_0_n_10), .D(watchdog_0_n_12), .RN(watchdog_0_n_29));
  INV_X1_LVT watchdog_0_i_24_0 (.ZN(watchdog_0_wdtcnt_nxt[0]), .A(
      watchdog_0_wdtcnt[0]));
  AND2_X1_LVT watchdog_0_i_21_1 (.ZN(watchdog_0_n_11), .A1(watchdog_0_n_21_0), 
      .A2(watchdog_0_wdtcnt_nxt[0]));
  DFFR_X1_LVT \watchdog_0_wdtcnt_reg[0] (.Q(watchdog_0_wdtcnt[0]), .QN(), .CK(
      watchdog_0_n_10), .D(watchdog_0_n_11), .RN(watchdog_0_n_29));
  HA_X1_LVT watchdog_0_i_24_1 (.CO(watchdog_0_n_24_0), .S(
      watchdog_0_wdtcnt_nxt[1]), .A(watchdog_0_wdtcnt[1]), .B(
      watchdog_0_wdtcnt[0]));
  HA_X1_LVT watchdog_0_i_24_2 (.CO(watchdog_0_n_24_1), .S(
      watchdog_0_wdtcnt_nxt[2]), .A(watchdog_0_wdtcnt[2]), .B(watchdog_0_n_24_0));
  HA_X1_LVT watchdog_0_i_24_3 (.CO(watchdog_0_n_24_2), .S(
      watchdog_0_wdtcnt_nxt[3]), .A(watchdog_0_wdtcnt[3]), .B(watchdog_0_n_24_1));
  HA_X1_LVT watchdog_0_i_24_4 (.CO(watchdog_0_n_24_3), .S(
      watchdog_0_wdtcnt_nxt[4]), .A(watchdog_0_wdtcnt[4]), .B(watchdog_0_n_24_2));
  HA_X1_LVT watchdog_0_i_24_5 (.CO(watchdog_0_n_24_4), .S(
      watchdog_0_wdtcnt_nxt[5]), .A(watchdog_0_wdtcnt[5]), .B(watchdog_0_n_24_3));
  HA_X1_LVT watchdog_0_i_24_6 (.CO(watchdog_0_n_24_5), .S(
      watchdog_0_wdtcnt_nxt[6]), .A(watchdog_0_wdtcnt[6]), .B(watchdog_0_n_24_4));
  INV_X1_LVT watchdog_0_i_28_4 (.ZN(watchdog_0_n_28_4), .A(
      watchdog_0_wdtcnt_nxt[6]));
  OR4_X1_LVT watchdog_0_i_28_5 (.ZN(watchdog_0_n_28_5), .A1(watchdog_0_n_28_1), 
      .A2(watchdog_0_n_28_2), .A3(watchdog_0_n_28_3), .A4(watchdog_0_n_28_4));
  AND2_X1_LVT watchdog_0_i_21_16 (.ZN(watchdog_0_n_26), .A1(watchdog_0_n_21_0), 
      .A2(watchdog_0_wdtcnt_nxt[15]));
  DFFR_X1_LVT \watchdog_0_wdtcnt_reg[15] (.Q(watchdog_0_wdtcnt[15]), .QN(), .CK(
      watchdog_0_n_10), .D(watchdog_0_n_26), .RN(watchdog_0_n_29));
  AND2_X1_LVT watchdog_0_i_21_15 (.ZN(watchdog_0_n_25), .A1(watchdog_0_n_21_0), 
      .A2(watchdog_0_wdtcnt_nxt[14]));
  DFFR_X1_LVT \watchdog_0_wdtcnt_reg[14] (.Q(watchdog_0_wdtcnt[14]), .QN(), .CK(
      watchdog_0_n_10), .D(watchdog_0_n_25), .RN(watchdog_0_n_29));
  AND2_X1_LVT watchdog_0_i_21_14 (.ZN(watchdog_0_n_24), .A1(watchdog_0_n_21_0), 
      .A2(watchdog_0_wdtcnt_nxt[13]));
  DFFR_X1_LVT \watchdog_0_wdtcnt_reg[13] (.Q(watchdog_0_wdtcnt[13]), .QN(), .CK(
      watchdog_0_n_10), .D(watchdog_0_n_24), .RN(watchdog_0_n_29));
  AND2_X1_LVT watchdog_0_i_21_13 (.ZN(watchdog_0_n_23), .A1(watchdog_0_n_21_0), 
      .A2(watchdog_0_wdtcnt_nxt[12]));
  DFFR_X1_LVT \watchdog_0_wdtcnt_reg[12] (.Q(watchdog_0_wdtcnt[12]), .QN(), .CK(
      watchdog_0_n_10), .D(watchdog_0_n_23), .RN(watchdog_0_n_29));
  AND2_X1_LVT watchdog_0_i_21_12 (.ZN(watchdog_0_n_22), .A1(watchdog_0_n_21_0), 
      .A2(watchdog_0_wdtcnt_nxt[11]));
  DFFR_X1_LVT \watchdog_0_wdtcnt_reg[11] (.Q(watchdog_0_wdtcnt[11]), .QN(), .CK(
      watchdog_0_n_10), .D(watchdog_0_n_22), .RN(watchdog_0_n_29));
  AND2_X1_LVT watchdog_0_i_21_11 (.ZN(watchdog_0_n_21), .A1(watchdog_0_n_21_0), 
      .A2(watchdog_0_wdtcnt_nxt[10]));
  DFFR_X1_LVT \watchdog_0_wdtcnt_reg[10] (.Q(watchdog_0_wdtcnt[10]), .QN(), .CK(
      watchdog_0_n_10), .D(watchdog_0_n_21), .RN(watchdog_0_n_29));
  AND2_X1_LVT watchdog_0_i_21_10 (.ZN(watchdog_0_n_20), .A1(watchdog_0_n_21_0), 
      .A2(watchdog_0_wdtcnt_nxt[9]));
  DFFR_X1_LVT \watchdog_0_wdtcnt_reg[9] (.Q(watchdog_0_wdtcnt[9]), .QN(), .CK(
      watchdog_0_n_10), .D(watchdog_0_n_20), .RN(watchdog_0_n_29));
  AND2_X1_LVT watchdog_0_i_21_9 (.ZN(watchdog_0_n_19), .A1(watchdog_0_n_21_0), 
      .A2(watchdog_0_wdtcnt_nxt[8]));
  DFFR_X1_LVT \watchdog_0_wdtcnt_reg[8] (.Q(watchdog_0_wdtcnt[8]), .QN(), .CK(
      watchdog_0_n_10), .D(watchdog_0_n_19), .RN(watchdog_0_n_29));
  AND2_X1_LVT watchdog_0_i_21_8 (.ZN(watchdog_0_n_18), .A1(watchdog_0_n_21_0), 
      .A2(watchdog_0_wdtcnt_nxt[7]));
  DFFR_X1_LVT \watchdog_0_wdtcnt_reg[7] (.Q(watchdog_0_wdtcnt[7]), .QN(), .CK(
      watchdog_0_n_10), .D(watchdog_0_n_18), .RN(watchdog_0_n_29));
  HA_X1_LVT watchdog_0_i_24_7 (.CO(watchdog_0_n_24_6), .S(
      watchdog_0_wdtcnt_nxt[7]), .A(watchdog_0_wdtcnt[7]), .B(watchdog_0_n_24_5));
  HA_X1_LVT watchdog_0_i_24_8 (.CO(watchdog_0_n_24_7), .S(
      watchdog_0_wdtcnt_nxt[8]), .A(watchdog_0_wdtcnt[8]), .B(watchdog_0_n_24_6));
  HA_X1_LVT watchdog_0_i_24_9 (.CO(watchdog_0_n_24_8), .S(
      watchdog_0_wdtcnt_nxt[9]), .A(watchdog_0_wdtcnt[9]), .B(watchdog_0_n_24_7));
  HA_X1_LVT watchdog_0_i_24_10 (.CO(watchdog_0_n_24_9), .S(
      watchdog_0_wdtcnt_nxt[10]), .A(watchdog_0_wdtcnt[10]), .B(
      watchdog_0_n_24_8));
  HA_X1_LVT watchdog_0_i_24_11 (.CO(watchdog_0_n_24_10), .S(
      watchdog_0_wdtcnt_nxt[11]), .A(watchdog_0_wdtcnt[11]), .B(
      watchdog_0_n_24_9));
  HA_X1_LVT watchdog_0_i_24_12 (.CO(watchdog_0_n_24_11), .S(
      watchdog_0_wdtcnt_nxt[12]), .A(watchdog_0_wdtcnt[12]), .B(
      watchdog_0_n_24_10));
  HA_X1_LVT watchdog_0_i_24_13 (.CO(watchdog_0_n_24_12), .S(
      watchdog_0_wdtcnt_nxt[13]), .A(watchdog_0_wdtcnt[13]), .B(
      watchdog_0_n_24_11));
  HA_X1_LVT watchdog_0_i_24_14 (.CO(watchdog_0_n_24_13), .S(
      watchdog_0_wdtcnt_nxt[14]), .A(watchdog_0_wdtcnt[14]), .B(
      watchdog_0_n_24_12));
  XNOR2_X1_LVT watchdog_0_i_24_15 (.ZN(watchdog_0_n_24_14), .A(
      watchdog_0_wdtcnt[15]), .B(watchdog_0_n_24_13));
  INV_X1_LVT watchdog_0_i_24_16 (.ZN(watchdog_0_wdtcnt_nxt[15]), .A(
      watchdog_0_n_24_14));
  NAND2_X1_LVT watchdog_0_i_28_6 (.ZN(watchdog_0_n_28_6), .A1(watchdog_0_n_28_3), 
      .A2(watchdog_0_wdtcnt_nxt[15]));
  NAND2_X1_LVT watchdog_0_i_28_7 (.ZN(watchdog_0_n_28_7), .A1(watchdog_0_n_28_2), 
      .A2(watchdog_0_wdtcnt_nxt[13]));
  NAND2_X1_LVT watchdog_0_i_28_8 (.ZN(watchdog_0_n_28_8), .A1(watchdog_0_n_28_1), 
      .A2(watchdog_0_wdtcnt_nxt[9]));
  NAND4_X1_LVT watchdog_0_i_28_9 (.ZN(watchdog_0_wdtqn_reg), .A1(
      watchdog_0_n_28_5), .A2(watchdog_0_n_28_6), .A3(watchdog_0_n_28_7), .A4(
      watchdog_0_n_28_8));
  AND2_X1_LVT watchdog_0_i_29_0 (.ZN(watchdog_0_wdtqn_edge), .A1(
      watchdog_0_wdtqn_reg), .A2(watchdog_0_wdtcnt_incr));
  CLKGATETST_X1_LVT watchdog_0_clk_gate_wdt_evt_toggle_reg (.GCK(watchdog_0_n_28), 
      .CK(smclk), .E(watchdog_0_wdtqn_edge), .SE(1'b0));
  DFFR_X1_LVT watchdog_0_wdt_evt_toggle_reg (.Q(watchdog_0_wdt_evt_toggle), .QN(), 
      .CK(watchdog_0_n_28), .D(watchdog_0_n_30), .RN(watchdog_0_n_29));
  INV_X1_LVT watchdog_0_sync_cell_wdt_evt_i_0_0 (.ZN(
      watchdog_0_sync_cell_wdt_evt_n_0), .A(puc_rst));
  DFFR_X1_LVT \watchdog_0_sync_cell_wdt_evt_data_sync_reg[0] (.Q(
      watchdog_0_sync_cell_wdt_evt_n_1), .QN(), .CK(mclk), .D(
      watchdog_0_wdt_evt_toggle), .RN(watchdog_0_sync_cell_wdt_evt_n_0));
  DFFR_X1_LVT \watchdog_0_sync_cell_wdt_evt_data_sync_reg[1] (.Q(
      watchdog_0_wdt_evt_toggle_sync), .QN(), .CK(mclk), .D(
      watchdog_0_sync_cell_wdt_evt_n_1), .RN(watchdog_0_sync_cell_wdt_evt_n_0));
  DFFR_X1_LVT watchdog_0_wdt_evt_toggle_sync_dly_reg (.Q(
      watchdog_0_wdt_evt_toggle_sync_dly), .QN(), .CK(mclk), .D(
      watchdog_0_wdt_evt_toggle_sync), .RN(watchdog_0_n_4));
  XOR2_X1_LVT watchdog_0_i_9_0 (.Z(watchdog_0_n_9_0), .A(
      watchdog_0_wdt_evt_toggle_sync_dly), .B(watchdog_0_wdt_evt_toggle_sync));
  INV_X1_LVT watchdog_0_i_8_0 (.ZN(watchdog_0_n_8_0), .A(watchdog_0_reg_wr));
  AND4_X1_LVT watchdog_0_i_8_1 (.ZN(watchdog_0_n_8_1), .A1(per_din[9]), .A2(
      per_din[11]), .A3(per_din[12]), .A4(per_din[14]));
  NOR4_X1_LVT watchdog_0_i_8_2 (.ZN(watchdog_0_n_8_2), .A1(per_din[8]), .A2(
      per_din[10]), .A3(per_din[13]), .A4(per_din[15]));
  AOI21_X1_LVT watchdog_0_i_8_3 (.ZN(watchdog_0_wdtpw_error), .A(
      watchdog_0_n_8_0), .B1(watchdog_0_n_8_1), .B2(watchdog_0_n_8_2));
  OR3_X1_LVT watchdog_0_i_9_1 (.ZN(watchdog_0_wdtifg_set), .A1(watchdog_0_n_9_0), 
      .A2(wdtifg_sw_set), .A3(watchdog_0_wdtpw_error));
  AOI21_X1_LVT watchdog_0_i_10_0 (.ZN(watchdog_0_n_10_0), .A(wdtifg_sw_clr), .B1(
      irq_acc[10]), .B2(watchdog_0_wdtctl[4]));
  INV_X1_LVT watchdog_0_i_10_1 (.ZN(watchdog_0_wdtifg_clr), .A(watchdog_0_n_10_0));
  INV_X1_LVT watchdog_0_i_13_1 (.ZN(watchdog_0_n_13_1), .A(watchdog_0_wdtifg_clr));
  INV_X1_LVT watchdog_0_i_13_0 (.ZN(watchdog_0_n_13_0), .A(watchdog_0_wdtifg_set));
  NAND2_X1_LVT watchdog_0_i_13_2 (.ZN(watchdog_0_n_7), .A1(watchdog_0_n_13_1), 
      .A2(watchdog_0_n_13_0));
  CLKGATETST_X1_LVT watchdog_0_clk_gate_wdtifg_reg (.GCK(watchdog_0_n_5), .CK(
      mclk), .E(watchdog_0_n_7), .SE(1'b0));
  INV_X1_LVT watchdog_0_i_11_0 (.ZN(watchdog_0_n_6), .A(por));
  DFFR_X1_LVT watchdog_0_wdtifg_reg (.Q(wdtifg), .QN(), .CK(watchdog_0_n_5), .D(
      watchdog_0_wdtifg_set), .RN(watchdog_0_n_6));
  AND3_X1_LVT watchdog_0_i_15_0 (.ZN(wdt_irq), .A1(watchdog_0_wdtctl[4]), .A2(
      wdtie), .A3(wdtifg));
  INV_X1_LVT watchdog_0_i_16_0 (.ZN(watchdog_0_n_8), .A(watchdog_0_wdtctl[4]));
  AOI21_X1_LVT watchdog_0_i_17_0 (.ZN(watchdog_0_n_17_0), .A(
      watchdog_0_wdtpw_error), .B1(watchdog_0_wdtifg_set), .B2(watchdog_0_n_8));
  INV_X1_LVT watchdog_0_i_17_1 (.ZN(watchdog_0_n_9), .A(watchdog_0_n_17_0));
  DFFR_X1_LVT watchdog_0_wdt_reset_reg (.Q(wdt_reset), .QN(), .CK(mclk), .D(
      watchdog_0_n_9), .RN(watchdog_0_n_6));
  DFFS_X1_LVT watchdog_0_wdtifg_clr_reg_reg (.Q(watchdog_0_wdtifg_clr_reg), .QN(), 
      .CK(mclk), .D(watchdog_0_wdtifg_clr), .SN(watchdog_0_n_4));
  DFFR_X1_LVT watchdog_0_wdtqn_edge_reg_reg (.Q(watchdog_0_wdtqn_edge_reg), .QN(), 
      .CK(smclk), .D(watchdog_0_wdtqn_edge), .RN(watchdog_0_n_29));
  INV_X1_LVT watchdog_0_wakeup_cell_wdog_scan_mux_clk_i_0_0 (.ZN(
      watchdog_0_wakeup_cell_wdog_scan_mux_clk_n_0_0), .A(scan_mode));
  AOI22_X1_LVT watchdog_0_wakeup_cell_wdog_scan_mux_clk_i_0_1 (.ZN(
      watchdog_0_wakeup_cell_wdog_scan_mux_clk_n_0_1), .A1(
      watchdog_0_wakeup_cell_wdog_scan_mux_clk_n_0_0), .A2(
      watchdog_0_wdtqn_edge_reg), .B1(mclk), .B2(scan_mode));
  INV_X1_LVT watchdog_0_wakeup_cell_wdog_scan_mux_clk_i_0_2 (.ZN(
      watchdog_0_wakeup_cell_wdog_wkup_clk), .A(
      watchdog_0_wakeup_cell_wdog_scan_mux_clk_n_0_1));
  INV_X1_LVT watchdog_0_wakeup_cell_wdog_scan_mux_rst_i_0_0 (.ZN(
      watchdog_0_wakeup_cell_wdog_scan_mux_rst_n_0_0), .A(scan_mode));
  AOI22_X1_LVT watchdog_0_wakeup_cell_wdog_scan_mux_rst_i_0_1 (.ZN(
      watchdog_0_wakeup_cell_wdog_scan_mux_rst_n_0_1), .A1(
      watchdog_0_wakeup_cell_wdog_scan_mux_rst_n_0_0), .A2(
      watchdog_0_wdtifg_clr_reg), .B1(puc_rst), .B2(scan_mode));
  INV_X1_LVT watchdog_0_wakeup_cell_wdog_scan_mux_rst_i_0_2 (.ZN(
      watchdog_0_wakeup_cell_wdog_wkup_rst), .A(
      watchdog_0_wakeup_cell_wdog_scan_mux_rst_n_0_1));
  INV_X1_LVT watchdog_0_wakeup_cell_wdog_i_0_0 (.ZN(
      watchdog_0_wakeup_cell_wdog_n_0), .A(watchdog_0_wakeup_cell_wdog_wkup_rst));
  DFFR_X1_LVT watchdog_0_wakeup_cell_wdog_wkup_out_reg (.Q(
      watchdog_0_wdt_wkup_pre), .QN(), .CK(watchdog_0_wakeup_cell_wdog_wkup_clk), 
      .D(1'b1), .RN(watchdog_0_wakeup_cell_wdog_n_0));
  NOR2_X1_LVT watchdog_0_i_35_2 (.ZN(watchdog_0_n_35_1), .A1(wdtie), .A2(
      watchdog_0_n_8));
  INV_X1_LVT watchdog_0_i_35_0 (.ZN(watchdog_0_n_35_0), .A(watchdog_0_n_31));
  NOR2_X1_LVT watchdog_0_i_35_1 (.ZN(watchdog_0_n_32), .A1(watchdog_0_n_35_1), 
      .A2(watchdog_0_n_35_0));
  DFFR_X1_LVT watchdog_0_wdt_wkup_en_reg (.Q(watchdog_0_wdt_wkup_en), .QN(), .CK(
      mclk), .D(watchdog_0_n_32), .RN(watchdog_0_n_4));
  AND2_X1_LVT watchdog_0_and_wdt_wkup_i_0_0 (.ZN(wdt_wkup), .A1(
      watchdog_0_wdt_wkup_pre), .A2(watchdog_0_wdt_wkup_en));
  DFFR_X1_LVT \watchdog_0_wdtctl_reg[5] (.Q(watchdog_0_wdtctl[5]), .QN(), .CK(
      watchdog_0_n_3), .D(1'b0), .RN(watchdog_0_n_4));
  INV_X1_LVT sfr_0_i_13_1 (.ZN(sfr_0_n_13_1), .A(per_din[4]));
  INV_X1_LVT sfr_0_i_0_0 (.ZN(sfr_0_n_0_0), .A(per_en));
  NOR4_X1_LVT sfr_0_i_0_1 (.ZN(sfr_0_n_0_1), .A1(sfr_0_n_0_0), .A2(per_addr[11]), 
      .A3(per_addr[12]), .A4(per_addr[13]));
  NOR4_X1_LVT sfr_0_i_0_2 (.ZN(sfr_0_n_0_2), .A1(per_addr[3]), .A2(per_addr[4]), 
      .A3(per_addr[5]), .A4(per_addr[6]));
  NOR4_X1_LVT sfr_0_i_0_3 (.ZN(sfr_0_n_0_3), .A1(per_addr[7]), .A2(per_addr[8]), 
      .A3(per_addr[9]), .A4(per_addr[10]));
  AND3_X1_LVT sfr_0_i_0_4 (.ZN(sfr_0_reg_sel), .A1(sfr_0_n_0_1), .A2(sfr_0_n_0_2), 
      .A3(sfr_0_n_0_3));
  AND2_X1_LVT sfr_0_i_1_0 (.ZN(sfr_0_reg_lo_write), .A1(per_we[0]), .A2(
      sfr_0_reg_sel));
  INV_X1_LVT sfr_0_i_2_1 (.ZN(sfr_0_n_2_1), .A(per_addr[1]));
  NAND2_X1_LVT sfr_0_i_2_3 (.ZN(sfr_0_n_2_3), .A1(per_addr[0]), .A2(sfr_0_n_2_1));
  NOR2_X1_LVT sfr_0_i_2_8 (.ZN(sfr_0_n_1), .A1(sfr_0_n_2_3), .A2(per_addr[2]));
  AND2_X1_LVT sfr_0_i_3_1 (.ZN(sfr_0_ifg1_wr), .A1(sfr_0_reg_lo_write), .A2(
      sfr_0_n_1));
  INV_X1_LVT sfr_0_i_4_0 (.ZN(sfr_0_n_4_0), .A(sfr_0_ifg1_wr));
  NOR2_X1_LVT sfr_0_i_4_1 (.ZN(sfr_0_n_6), .A1(sfr_0_n_4_0), .A2(per_din[4]));
  INV_X1_LVT sfr_0_i_11_0 (.ZN(sfr_0_n_11), .A(puc_rst));
  DFFS_X1_LVT sfr_0_nmi_capture_rst_reg (.Q(sfr_0_nmi_capture_rst), .QN(), .CK(
      mclk), .D(sfr_0_n_6), .SN(sfr_0_n_11));
  XOR2_X1_LVT sfr_0_i_31_0 (.Z(sfr_0_nmi_pol), .A(nmi), .B(wdtnmies));
  INV_X1_LVT sfr_0_wakeup_cell_nmi_scan_mux_clk_i_0_0 (.ZN(
      sfr_0_wakeup_cell_nmi_scan_mux_clk_n_0_0), .A(scan_mode));
  AOI22_X1_LVT sfr_0_wakeup_cell_nmi_scan_mux_clk_i_0_1 (.ZN(
      sfr_0_wakeup_cell_nmi_scan_mux_clk_n_0_1), .A1(
      sfr_0_wakeup_cell_nmi_scan_mux_clk_n_0_0), .A2(sfr_0_nmi_pol), .B1(mclk), 
      .B2(scan_mode));
  INV_X1_LVT sfr_0_wakeup_cell_nmi_scan_mux_clk_i_0_2 (.ZN(
      sfr_0_wakeup_cell_nmi_wkup_clk), .A(
      sfr_0_wakeup_cell_nmi_scan_mux_clk_n_0_1));
  INV_X1_LVT sfr_0_wakeup_cell_nmi_scan_mux_rst_i_0_0 (.ZN(
      sfr_0_wakeup_cell_nmi_scan_mux_rst_n_0_0), .A(scan_mode));
  AOI22_X1_LVT sfr_0_wakeup_cell_nmi_scan_mux_rst_i_0_1 (.ZN(
      sfr_0_wakeup_cell_nmi_scan_mux_rst_n_0_1), .A1(
      sfr_0_wakeup_cell_nmi_scan_mux_rst_n_0_0), .A2(sfr_0_nmi_capture_rst), .B1(
      puc_rst), .B2(scan_mode));
  INV_X1_LVT sfr_0_wakeup_cell_nmi_scan_mux_rst_i_0_2 (.ZN(
      sfr_0_wakeup_cell_nmi_wkup_rst), .A(
      sfr_0_wakeup_cell_nmi_scan_mux_rst_n_0_1));
  INV_X1_LVT sfr_0_wakeup_cell_nmi_i_0_0 (.ZN(sfr_0_wakeup_cell_nmi_n_0), .A(
      sfr_0_wakeup_cell_nmi_wkup_rst));
  DFFR_X1_LVT sfr_0_wakeup_cell_nmi_wkup_out_reg (.Q(sfr_0_nmi_capture), .QN(), 
      .CK(sfr_0_wakeup_cell_nmi_wkup_clk), .D(1'b1), .RN(
      sfr_0_wakeup_cell_nmi_n_0));
  INV_X1_LVT sfr_0_sync_cell_nmi_i_0_0 (.ZN(sfr_0_sync_cell_nmi_n_0), .A(puc_rst));
  DFFR_X1_LVT \sfr_0_sync_cell_nmi_data_sync_reg[0] (.Q(sfr_0_sync_cell_nmi_n_1), 
      .QN(), .CK(mclk), .D(sfr_0_nmi_capture), .RN(sfr_0_sync_cell_nmi_n_0));
  DFFR_X1_LVT \sfr_0_sync_cell_nmi_data_sync_reg[1] (.Q(sfr_0_nmi_s), .QN(), .CK(
      mclk), .D(sfr_0_sync_cell_nmi_n_1), .RN(sfr_0_sync_cell_nmi_n_0));
  INV_X1_LVT sfr_0_i_10_0 (.ZN(sfr_0_n_10_0), .A(sfr_0_nmi_s));
  DFFR_X1_LVT sfr_0_nmi_dly_reg (.Q(sfr_0_nmi_dly), .QN(), .CK(mclk), .D(
      sfr_0_nmi_s), .RN(sfr_0_n_11));
  NOR2_X1_LVT sfr_0_i_10_1 (.ZN(sfr_0_nmi_edge), .A1(sfr_0_n_10_0), .A2(
      sfr_0_nmi_dly));
  INV_X1_LVT sfr_0_i_13_0 (.ZN(sfr_0_n_13_0), .A(sfr_0_nmi_edge));
  NAND2_X1_LVT sfr_0_i_13_2 (.ZN(sfr_0_n_12), .A1(sfr_0_n_13_1), .A2(
      sfr_0_n_13_0));
  INV_X1_LVT sfr_0_i_14_1 (.ZN(sfr_0_n_14_1), .A(sfr_0_ifg1_wr));
  INV_X1_LVT sfr_0_i_14_0 (.ZN(sfr_0_n_14_0), .A(sfr_0_nmi_edge));
  NAND2_X1_LVT sfr_0_i_14_2 (.ZN(sfr_0_n_13), .A1(sfr_0_n_14_1), .A2(
      sfr_0_n_14_0));
  CLKGATETST_X1_LVT sfr_0_clk_gate_nmiifg_reg (.GCK(sfr_0_n_10), .CK(mclk), .E(
      sfr_0_n_13), .SE(1'b0));
  DFFR_X1_LVT sfr_0_nmiifg_reg (.Q(sfr_0_nmiifg), .QN(), .CK(sfr_0_n_10), .D(
      sfr_0_n_12), .RN(sfr_0_n_11));
  INV_X1_LVT sfr_0_i_7_0 (.ZN(sfr_0_n_7_0), .A(per_din[4]));
  NOR2_X1_LVT sfr_0_i_7_1 (.ZN(sfr_0_n_8), .A1(sfr_0_n_7_0), .A2(nmi_acc));
  INV_X1_LVT sfr_0_i_2_0 (.ZN(sfr_0_n_2_0), .A(per_addr[0]));
  NAND2_X1_LVT sfr_0_i_2_2 (.ZN(sfr_0_n_2_2), .A1(sfr_0_n_2_0), .A2(sfr_0_n_2_1));
  NOR2_X1_LVT sfr_0_i_2_7 (.ZN(sfr_0_n_0), .A1(sfr_0_n_2_2), .A2(per_addr[2]));
  AND2_X1_LVT sfr_0_i_3_0 (.ZN(sfr_0_n_5), .A1(sfr_0_n_0), .A2(
      sfr_0_reg_lo_write));
  INV_X1_LVT sfr_0_i_8_1 (.ZN(sfr_0_n_8_1), .A(sfr_0_n_5));
  INV_X1_LVT sfr_0_i_8_0 (.ZN(sfr_0_n_8_0), .A(nmi_acc));
  NAND2_X1_LVT sfr_0_i_8_2 (.ZN(sfr_0_n_9), .A1(sfr_0_n_8_1), .A2(sfr_0_n_8_0));
  CLKGATETST_X1_LVT sfr_0_clk_gate_nmie_reg (.GCK(sfr_0_n_7), .CK(mclk), .E(
      sfr_0_n_9), .SE(1'b0));
  DFFR_X1_LVT sfr_0_nmie_reg (.Q(sfr_0_nmie), .QN(), .CK(sfr_0_n_7), .D(
      sfr_0_n_8), .RN(sfr_0_n_11));
  AND2_X1_LVT sfr_0_i_16_0 (.ZN(nmi_pnd), .A1(sfr_0_nmiifg), .A2(sfr_0_nmie));
  XOR2_X1_LVT sfr_0_i_30_0 (.Z(sfr_0_n_31), .A(sfr_0_nmi_capture), .B(
      sfr_0_nmi_dly));
  AND2_X1_LVT sfr_0_and_nmi_wkup_i_0_0 (.ZN(nmi_wkup), .A1(sfr_0_n_31), .A2(
      sfr_0_nmie));
  NOR2_X1_LVT sfr_0_i_17_0 (.ZN(sfr_0_n_14), .A1(per_we[0]), .A2(per_we[1]));
  AND2_X1_LVT sfr_0_i_18_0 (.ZN(sfr_0_reg_read), .A1(sfr_0_n_14), .A2(
      sfr_0_reg_sel));
  INV_X1_LVT sfr_0_i_2_6 (.ZN(sfr_0_n_2_6), .A(per_addr[2]));
  NOR2_X1_LVT sfr_0_i_2_11 (.ZN(sfr_0_n_4), .A1(sfr_0_n_2_2), .A2(sfr_0_n_2_6));
  AND2_X1_LVT sfr_0_i_19_4 (.ZN(sfr_0_n_19), .A1(sfr_0_reg_read), .A2(sfr_0_n_4));
  AND2_X1_LVT sfr_0_i_21_7 (.ZN(per_dout_sfr[15]), .A1(sfr_0_n_19), .A2(1'b0));
  AND2_X1_LVT sfr_0_i_21_6 (.ZN(per_dout_sfr[14]), .A1(sfr_0_n_19), .A2(1'b0));
  AND2_X1_LVT sfr_0_i_21_5 (.ZN(per_dout_sfr[13]), .A1(sfr_0_n_19), .A2(1'b0));
  NAND2_X1_LVT sfr_0_i_2_5 (.ZN(sfr_0_n_2_5), .A1(per_addr[0]), .A2(per_addr[1]));
  NOR2_X1_LVT sfr_0_i_2_10 (.ZN(sfr_0_n_3), .A1(sfr_0_n_2_5), .A2(per_addr[2]));
  AND2_X1_LVT sfr_0_i_19_3 (.ZN(sfr_0_n_18), .A1(sfr_0_reg_read), .A2(sfr_0_n_3));
  AND2_X1_LVT sfr_0_i_21_4 (.ZN(sfr_0_n_25), .A1(sfr_0_n_19), .A2(1'b0));
  OR2_X1_LVT sfr_0_i_27_6 (.ZN(per_dout_sfr[12]), .A1(sfr_0_n_18), .A2(
      sfr_0_n_25));
  AND2_X1_LVT sfr_0_i_21_3 (.ZN(per_dout_sfr[11]), .A1(sfr_0_n_19), .A2(1'b0));
  AND2_X1_LVT sfr_0_i_21_2 (.ZN(per_dout_sfr[10]), .A1(sfr_0_n_19), .A2(1'b0));
  NAND2_X1_LVT sfr_0_i_2_4 (.ZN(sfr_0_n_2_4), .A1(sfr_0_n_2_0), .A2(per_addr[1]));
  NOR2_X1_LVT sfr_0_i_2_9 (.ZN(sfr_0_n_2), .A1(sfr_0_n_2_4), .A2(per_addr[2]));
  AND2_X1_LVT sfr_0_i_19_2 (.ZN(sfr_0_n_17), .A1(sfr_0_reg_read), .A2(sfr_0_n_2));
  AND2_X1_LVT sfr_0_i_21_1 (.ZN(sfr_0_n_24), .A1(sfr_0_n_19), .A2(1'b0));
  OR2_X1_LVT sfr_0_i_27_5 (.ZN(per_dout_sfr[9]), .A1(sfr_0_n_17), .A2(sfr_0_n_24));
  AND2_X1_LVT sfr_0_i_21_0 (.ZN(per_dout_sfr[8]), .A1(1'b0), .A2(sfr_0_n_19));
  AND2_X1_LVT sfr_0_i_20_7 (.ZN(per_dout_sfr[7]), .A1(sfr_0_n_19), .A2(1'b0));
  AND2_X1_LVT sfr_0_i_20_6 (.ZN(per_dout_sfr[6]), .A1(sfr_0_n_19), .A2(1'b0));
  AND2_X1_LVT sfr_0_i_20_5 (.ZN(per_dout_sfr[5]), .A1(sfr_0_n_19), .A2(1'b0));
  AND2_X1_LVT sfr_0_i_19_0 (.ZN(sfr_0_n_15), .A1(sfr_0_n_0), .A2(sfr_0_reg_read));
  AND2_X1_LVT sfr_0_i_26_0 (.ZN(sfr_0_n_30), .A1(sfr_0_nmie), .A2(sfr_0_n_15));
  AND2_X1_LVT sfr_0_i_19_1 (.ZN(sfr_0_n_16), .A1(sfr_0_reg_read), .A2(sfr_0_n_1));
  AND2_X1_LVT sfr_0_i_23_0 (.ZN(sfr_0_n_27), .A1(sfr_0_nmiifg), .A2(sfr_0_n_16));
  AND2_X1_LVT sfr_0_i_20_4 (.ZN(sfr_0_n_23), .A1(sfr_0_n_19), .A2(1'b0));
  OR4_X1_LVT sfr_0_i_27_4 (.ZN(per_dout_sfr[4]), .A1(sfr_0_n_30), .A2(sfr_0_n_27), 
      .A3(sfr_0_n_18), .A4(sfr_0_n_23));
  AND2_X1_LVT sfr_0_i_20_3 (.ZN(sfr_0_n_22), .A1(sfr_0_n_19), .A2(1'b0));
  OR2_X1_LVT sfr_0_i_27_3 (.ZN(per_dout_sfr[3]), .A1(sfr_0_n_17), .A2(sfr_0_n_22));
  AND2_X1_LVT sfr_0_i_20_2 (.ZN(per_dout_sfr[2]), .A1(sfr_0_n_19), .A2(1'b0));
  AND2_X1_LVT sfr_0_i_20_1 (.ZN(sfr_0_n_21), .A1(sfr_0_n_19), .A2(1'b0));
  OR2_X1_LVT sfr_0_i_27_2 (.ZN(per_dout_sfr[1]), .A1(sfr_0_n_17), .A2(sfr_0_n_21));
  AND2_X1_LVT sfr_0_i_22_0 (.ZN(sfr_0_n_26), .A1(wdtifg), .A2(sfr_0_n_16));
  AND2_X1_LVT sfr_0_i_20_0 (.ZN(sfr_0_n_20), .A1(1'b0), .A2(sfr_0_n_19));
  OR4_X1_LVT sfr_0_i_27_0 (.ZN(sfr_0_n_27_0), .A1(sfr_0_n_26), .A2(sfr_0_n_17), 
      .A3(sfr_0_n_18), .A4(sfr_0_n_20));
  CLKGATETST_X1_LVT sfr_0_clk_gate_wdtie_reg (.GCK(sfr_0_n_28), .CK(mclk), .E(
      sfr_0_n_5), .SE(1'b0));
  DFFR_X1_LVT sfr_0_wdtie_reg (.Q(wdtie), .QN(), .CK(sfr_0_n_28), .D(per_din[0]), 
      .RN(sfr_0_n_11));
  AND2_X1_LVT sfr_0_i_25_0 (.ZN(sfr_0_n_29), .A1(wdtie), .A2(sfr_0_n_15));
  OR2_X1_LVT sfr_0_i_27_1 (.ZN(per_dout_sfr[0]), .A1(sfr_0_n_27_0), .A2(
      sfr_0_n_29));
  INV_X1_LVT sfr_0_i_28_0 (.ZN(sfr_0_n_28_0), .A(sfr_0_ifg1_wr));
  NOR2_X1_LVT sfr_0_i_28_1 (.ZN(wdtifg_sw_clr), .A1(sfr_0_n_28_0), .A2(per_din[0]));
  AND2_X1_LVT sfr_0_i_29_0 (.ZN(wdtifg_sw_set), .A1(sfr_0_ifg1_wr), .A2(
      per_din[0]));
  INV_X1_LVT dbg_0_i_48_2 (.ZN(dbg_0_n_48_1), .A(dbg_0_dbg_addr[1]));
  NAND2_X1_LVT dbg_0_i_48_7 (.ZN(dbg_0_dbg_addr_in[1]), .A1(dbg_0_n_48_1), .A2(
      dbg_0_n_48_0));
  NOR2_X1_LVT dbg_0_i_49_2 (.ZN(dbg_0_n_49_2), .A1(dbg_0_dbg_addr_in[0]), .A2(
      dbg_0_dbg_addr_in[1]));
  INV_X1_LVT dbg_0_i_48_3 (.ZN(dbg_0_n_48_2), .A(dbg_0_dbg_addr[2]));
  NAND2_X1_LVT dbg_0_i_48_8 (.ZN(dbg_0_dbg_addr_in[2]), .A1(dbg_0_n_48_2), .A2(
      dbg_0_n_48_0));
  NAND2_X1_LVT dbg_0_i_49_11 (.ZN(dbg_0_n_49_11), .A1(dbg_0_n_49_2), .A2(
      dbg_0_dbg_addr_in[2]));
  AND2_X1_LVT dbg_0_i_48_4 (.ZN(dbg_0_dbg_addr_in[3]), .A1(dbg_0_n_48_0), .A2(
      dbg_0_dbg_addr[3]));
  INV_X1_LVT dbg_0_i_49_15 (.ZN(dbg_0_n_49_15), .A(dbg_0_dbg_addr_in[3]));
  AND2_X1_LVT dbg_0_i_48_5 (.ZN(dbg_0_dbg_addr_in[4]), .A1(dbg_0_n_48_0), .A2(
      dbg_0_dbg_addr[4]));
  AND2_X1_LVT dbg_0_i_48_6 (.ZN(dbg_0_dbg_addr_in[5]), .A1(dbg_0_n_48_0), .A2(
      dbg_0_dbg_addr[5]));
  NOR2_X1_LVT dbg_0_i_49_16 (.ZN(dbg_0_n_49_16), .A1(dbg_0_dbg_addr_in[4]), .A2(
      dbg_0_dbg_addr_in[5]));
  NAND2_X1_LVT dbg_0_i_49_20 (.ZN(dbg_0_n_49_20), .A1(dbg_0_n_49_15), .A2(
      dbg_0_n_49_16));
  NOR2_X1_LVT dbg_0_i_49_26 (.ZN(dbg_0_n_95), .A1(dbg_0_n_49_11), .A2(
      dbg_0_n_49_20));
  AND2_X1_LVT dbg_0_i_50_2 (.ZN(dbg_0_mem_ctl_wr), .A1(dbg_0_dbg_wr), .A2(
      dbg_0_n_95));
  AND2_X1_LVT dbg_0_i_1_0 (.ZN(dbg_0_n_1), .A1(dbg_0_mem_ctl_wr), .A2(
      dbg_0_dbg_din[0]));
  INV_X1_LVT dbg_0_i_51_0 (.ZN(dbg_0_n_104), .A(dbg_rst));
  DFFR_X1_LVT dbg_0_mem_start_reg (.Q(dbg_0_mem_start), .QN(), .CK(dbg_clk), .D(
      dbg_0_n_1), .RN(dbg_0_n_104));
  AND2_X1_LVT dbg_0_i_50_5 (.ZN(dbg_0_n_102), .A1(dbg_0_dbg_wr), .A2(dbg_0_n_98));
  INV_X1_LVT dbg_0_i_40_0 (.ZN(dbg_0_n_40_0), .A(dbg_0_n_102));
  INV_X1_LVT dbg_0_i_39_3 (.ZN(dbg_0_n_39_2), .A(dbg_0_mem_cnt[0]));
  NAND2_X1_LVT dbg_0_i_39_2 (.ZN(dbg_0_n_39_1), .A1(dbg_0_n_55), .A2(
      dbg_0_n_39_2));
  XNOR2_X1_LVT dbg_0_i_39_4 (.ZN(dbg_0_n_57), .A(dbg_0_mem_cnt[1]), .B(
      dbg_0_n_39_1));
  AOI22_X1_LVT dbg_0_i_40_3 (.ZN(dbg_0_n_40_2), .A1(dbg_0_n_40_0), .A2(
      dbg_0_n_57), .B1(dbg_0_n_102), .B2(dbg_0_dbg_din[1]));
  INV_X1_LVT dbg_0_i_40_4 (.ZN(dbg_0_n_73), .A(dbg_0_n_40_2));
  DFFR_X1_LVT \dbg_0_mem_cnt_reg[1] (.Q(dbg_0_mem_cnt[1]), .QN(), .CK(dbg_clk), 
      .D(dbg_0_n_73), .RN(dbg_0_n_104));
  OR2_X1_LVT dbg_0_i_39_5 (.ZN(dbg_0_n_39_3), .A1(dbg_0_mem_cnt[1]), .A2(
      dbg_0_n_39_1));
  XNOR2_X1_LVT dbg_0_i_39_6 (.ZN(dbg_0_n_58), .A(dbg_0_mem_cnt[2]), .B(
      dbg_0_n_39_3));
  AOI22_X1_LVT dbg_0_i_40_5 (.ZN(dbg_0_n_40_3), .A1(dbg_0_n_40_0), .A2(
      dbg_0_n_58), .B1(dbg_0_n_102), .B2(dbg_0_dbg_din[2]));
  INV_X1_LVT dbg_0_i_40_6 (.ZN(dbg_0_n_74), .A(dbg_0_n_40_3));
  DFFR_X1_LVT \dbg_0_mem_cnt_reg[2] (.Q(dbg_0_mem_cnt[2]), .QN(), .CK(dbg_clk), 
      .D(dbg_0_n_74), .RN(dbg_0_n_104));
  OR2_X1_LVT dbg_0_i_39_7 (.ZN(dbg_0_n_39_4), .A1(dbg_0_mem_cnt[2]), .A2(
      dbg_0_n_39_3));
  XNOR2_X1_LVT dbg_0_i_39_8 (.ZN(dbg_0_n_59), .A(dbg_0_mem_cnt[3]), .B(
      dbg_0_n_39_4));
  AOI22_X1_LVT dbg_0_i_40_7 (.ZN(dbg_0_n_40_4), .A1(dbg_0_n_40_0), .A2(
      dbg_0_n_59), .B1(dbg_0_n_102), .B2(dbg_0_dbg_din[3]));
  INV_X1_LVT dbg_0_i_40_8 (.ZN(dbg_0_n_75), .A(dbg_0_n_40_4));
  DFFR_X1_LVT \dbg_0_mem_cnt_reg[3] (.Q(dbg_0_mem_cnt[3]), .QN(), .CK(dbg_clk), 
      .D(dbg_0_n_75), .RN(dbg_0_n_104));
  NOR4_X1_LVT dbg_0_i_37_0 (.ZN(dbg_0_n_37_0), .A1(dbg_0_mem_cnt[0]), .A2(
      dbg_0_mem_cnt[1]), .A3(dbg_0_mem_cnt[2]), .A4(dbg_0_mem_cnt[3]));
  OR2_X1_LVT dbg_0_i_39_9 (.ZN(dbg_0_n_39_5), .A1(dbg_0_mem_cnt[3]), .A2(
      dbg_0_n_39_4));
  XNOR2_X1_LVT dbg_0_i_39_10 (.ZN(dbg_0_n_60), .A(dbg_0_mem_cnt[4]), .B(
      dbg_0_n_39_5));
  AOI22_X1_LVT dbg_0_i_40_9 (.ZN(dbg_0_n_40_5), .A1(dbg_0_n_40_0), .A2(
      dbg_0_n_60), .B1(dbg_0_n_102), .B2(dbg_0_dbg_din[4]));
  INV_X1_LVT dbg_0_i_40_10 (.ZN(dbg_0_n_76), .A(dbg_0_n_40_5));
  DFFR_X1_LVT \dbg_0_mem_cnt_reg[4] (.Q(dbg_0_mem_cnt[4]), .QN(), .CK(dbg_clk), 
      .D(dbg_0_n_76), .RN(dbg_0_n_104));
  OR2_X1_LVT dbg_0_i_39_11 (.ZN(dbg_0_n_39_6), .A1(dbg_0_mem_cnt[4]), .A2(
      dbg_0_n_39_5));
  XNOR2_X1_LVT dbg_0_i_39_12 (.ZN(dbg_0_n_61), .A(dbg_0_mem_cnt[5]), .B(
      dbg_0_n_39_6));
  AOI22_X1_LVT dbg_0_i_40_11 (.ZN(dbg_0_n_40_6), .A1(dbg_0_n_40_0), .A2(
      dbg_0_n_61), .B1(dbg_0_n_102), .B2(dbg_0_dbg_din[5]));
  INV_X1_LVT dbg_0_i_40_12 (.ZN(dbg_0_n_77), .A(dbg_0_n_40_6));
  DFFR_X1_LVT \dbg_0_mem_cnt_reg[5] (.Q(dbg_0_mem_cnt[5]), .QN(), .CK(dbg_clk), 
      .D(dbg_0_n_77), .RN(dbg_0_n_104));
  OR2_X1_LVT dbg_0_i_39_13 (.ZN(dbg_0_n_39_7), .A1(dbg_0_mem_cnt[5]), .A2(
      dbg_0_n_39_6));
  XNOR2_X1_LVT dbg_0_i_39_14 (.ZN(dbg_0_n_62), .A(dbg_0_mem_cnt[6]), .B(
      dbg_0_n_39_7));
  AOI22_X1_LVT dbg_0_i_40_13 (.ZN(dbg_0_n_40_7), .A1(dbg_0_n_40_0), .A2(
      dbg_0_n_62), .B1(dbg_0_n_102), .B2(dbg_0_dbg_din[6]));
  INV_X1_LVT dbg_0_i_40_14 (.ZN(dbg_0_n_78), .A(dbg_0_n_40_7));
  DFFR_X1_LVT \dbg_0_mem_cnt_reg[6] (.Q(dbg_0_mem_cnt[6]), .QN(), .CK(dbg_clk), 
      .D(dbg_0_n_78), .RN(dbg_0_n_104));
  OR2_X1_LVT dbg_0_i_39_15 (.ZN(dbg_0_n_39_8), .A1(dbg_0_mem_cnt[6]), .A2(
      dbg_0_n_39_7));
  XNOR2_X1_LVT dbg_0_i_39_16 (.ZN(dbg_0_n_63), .A(dbg_0_mem_cnt[7]), .B(
      dbg_0_n_39_8));
  AOI22_X1_LVT dbg_0_i_40_15 (.ZN(dbg_0_n_40_8), .A1(dbg_0_n_40_0), .A2(
      dbg_0_n_63), .B1(dbg_0_n_102), .B2(dbg_0_dbg_din[7]));
  INV_X1_LVT dbg_0_i_40_16 (.ZN(dbg_0_n_79), .A(dbg_0_n_40_8));
  DFFR_X1_LVT \dbg_0_mem_cnt_reg[7] (.Q(dbg_0_mem_cnt[7]), .QN(), .CK(dbg_clk), 
      .D(dbg_0_n_79), .RN(dbg_0_n_104));
  NOR4_X1_LVT dbg_0_i_37_1 (.ZN(dbg_0_n_37_1), .A1(dbg_0_mem_cnt[4]), .A2(
      dbg_0_mem_cnt[5]), .A3(dbg_0_mem_cnt[6]), .A4(dbg_0_mem_cnt[7]));
  OR2_X1_LVT dbg_0_i_39_17 (.ZN(dbg_0_n_39_9), .A1(dbg_0_mem_cnt[7]), .A2(
      dbg_0_n_39_8));
  XNOR2_X1_LVT dbg_0_i_39_18 (.ZN(dbg_0_n_64), .A(dbg_0_mem_cnt[8]), .B(
      dbg_0_n_39_9));
  AOI22_X1_LVT dbg_0_i_40_17 (.ZN(dbg_0_n_40_9), .A1(dbg_0_n_40_0), .A2(
      dbg_0_n_64), .B1(dbg_0_n_102), .B2(dbg_0_dbg_din[8]));
  INV_X1_LVT dbg_0_i_40_18 (.ZN(dbg_0_n_80), .A(dbg_0_n_40_9));
  DFFR_X1_LVT \dbg_0_mem_cnt_reg[8] (.Q(dbg_0_mem_cnt[8]), .QN(), .CK(dbg_clk), 
      .D(dbg_0_n_80), .RN(dbg_0_n_104));
  OR2_X1_LVT dbg_0_i_39_19 (.ZN(dbg_0_n_39_10), .A1(dbg_0_mem_cnt[8]), .A2(
      dbg_0_n_39_9));
  XNOR2_X1_LVT dbg_0_i_39_20 (.ZN(dbg_0_n_65), .A(dbg_0_mem_cnt[9]), .B(
      dbg_0_n_39_10));
  AOI22_X1_LVT dbg_0_i_40_19 (.ZN(dbg_0_n_40_10), .A1(dbg_0_n_40_0), .A2(
      dbg_0_n_65), .B1(dbg_0_n_102), .B2(dbg_0_dbg_din[9]));
  INV_X1_LVT dbg_0_i_40_20 (.ZN(dbg_0_n_81), .A(dbg_0_n_40_10));
  DFFR_X1_LVT \dbg_0_mem_cnt_reg[9] (.Q(dbg_0_mem_cnt[9]), .QN(), .CK(dbg_clk), 
      .D(dbg_0_n_81), .RN(dbg_0_n_104));
  OR2_X1_LVT dbg_0_i_39_21 (.ZN(dbg_0_n_39_11), .A1(dbg_0_mem_cnt[9]), .A2(
      dbg_0_n_39_10));
  XNOR2_X1_LVT dbg_0_i_39_22 (.ZN(dbg_0_n_66), .A(dbg_0_mem_cnt[10]), .B(
      dbg_0_n_39_11));
  AOI22_X1_LVT dbg_0_i_40_21 (.ZN(dbg_0_n_40_11), .A1(dbg_0_n_40_0), .A2(
      dbg_0_n_66), .B1(dbg_0_n_102), .B2(dbg_0_dbg_din[10]));
  INV_X1_LVT dbg_0_i_40_22 (.ZN(dbg_0_n_82), .A(dbg_0_n_40_11));
  DFFR_X1_LVT \dbg_0_mem_cnt_reg[10] (.Q(dbg_0_mem_cnt[10]), .QN(), .CK(dbg_clk), 
      .D(dbg_0_n_82), .RN(dbg_0_n_104));
  OR2_X1_LVT dbg_0_i_39_23 (.ZN(dbg_0_n_39_12), .A1(dbg_0_mem_cnt[10]), .A2(
      dbg_0_n_39_11));
  XNOR2_X1_LVT dbg_0_i_39_24 (.ZN(dbg_0_n_67), .A(dbg_0_mem_cnt[11]), .B(
      dbg_0_n_39_12));
  AOI22_X1_LVT dbg_0_i_40_23 (.ZN(dbg_0_n_40_12), .A1(dbg_0_n_40_0), .A2(
      dbg_0_n_67), .B1(dbg_0_n_102), .B2(dbg_0_dbg_din[11]));
  INV_X1_LVT dbg_0_i_40_24 (.ZN(dbg_0_n_83), .A(dbg_0_n_40_12));
  DFFR_X1_LVT \dbg_0_mem_cnt_reg[11] (.Q(dbg_0_mem_cnt[11]), .QN(), .CK(dbg_clk), 
      .D(dbg_0_n_83), .RN(dbg_0_n_104));
  NOR4_X1_LVT dbg_0_i_37_2 (.ZN(dbg_0_n_37_2), .A1(dbg_0_mem_cnt[8]), .A2(
      dbg_0_mem_cnt[9]), .A3(dbg_0_mem_cnt[10]), .A4(dbg_0_mem_cnt[11]));
  OR2_X1_LVT dbg_0_i_39_25 (.ZN(dbg_0_n_39_13), .A1(dbg_0_mem_cnt[11]), .A2(
      dbg_0_n_39_12));
  XNOR2_X1_LVT dbg_0_i_39_26 (.ZN(dbg_0_n_68), .A(dbg_0_mem_cnt[12]), .B(
      dbg_0_n_39_13));
  AOI22_X1_LVT dbg_0_i_40_25 (.ZN(dbg_0_n_40_13), .A1(dbg_0_n_40_0), .A2(
      dbg_0_n_68), .B1(dbg_0_n_102), .B2(dbg_0_dbg_din[12]));
  INV_X1_LVT dbg_0_i_40_26 (.ZN(dbg_0_n_84), .A(dbg_0_n_40_13));
  DFFR_X1_LVT \dbg_0_mem_cnt_reg[12] (.Q(dbg_0_mem_cnt[12]), .QN(), .CK(dbg_clk), 
      .D(dbg_0_n_84), .RN(dbg_0_n_104));
  OR2_X1_LVT dbg_0_i_39_27 (.ZN(dbg_0_n_39_14), .A1(dbg_0_mem_cnt[12]), .A2(
      dbg_0_n_39_13));
  XNOR2_X1_LVT dbg_0_i_39_28 (.ZN(dbg_0_n_69), .A(dbg_0_mem_cnt[13]), .B(
      dbg_0_n_39_14));
  AOI22_X1_LVT dbg_0_i_40_27 (.ZN(dbg_0_n_40_14), .A1(dbg_0_n_40_0), .A2(
      dbg_0_n_69), .B1(dbg_0_n_102), .B2(dbg_0_dbg_din[13]));
  INV_X1_LVT dbg_0_i_40_28 (.ZN(dbg_0_n_85), .A(dbg_0_n_40_14));
  DFFR_X1_LVT \dbg_0_mem_cnt_reg[13] (.Q(dbg_0_mem_cnt[13]), .QN(), .CK(dbg_clk), 
      .D(dbg_0_n_85), .RN(dbg_0_n_104));
  OR2_X1_LVT dbg_0_i_39_29 (.ZN(dbg_0_n_39_15), .A1(dbg_0_mem_cnt[13]), .A2(
      dbg_0_n_39_14));
  XNOR2_X1_LVT dbg_0_i_39_30 (.ZN(dbg_0_n_70), .A(dbg_0_mem_cnt[14]), .B(
      dbg_0_n_39_15));
  AOI22_X1_LVT dbg_0_i_40_29 (.ZN(dbg_0_n_40_15), .A1(dbg_0_n_40_0), .A2(
      dbg_0_n_70), .B1(dbg_0_n_102), .B2(dbg_0_dbg_din[14]));
  INV_X1_LVT dbg_0_i_40_30 (.ZN(dbg_0_n_86), .A(dbg_0_n_40_15));
  DFFR_X1_LVT \dbg_0_mem_cnt_reg[14] (.Q(dbg_0_mem_cnt[14]), .QN(), .CK(dbg_clk), 
      .D(dbg_0_n_86), .RN(dbg_0_n_104));
  OR2_X1_LVT dbg_0_i_39_31 (.ZN(dbg_0_n_39_16), .A1(dbg_0_mem_cnt[14]), .A2(
      dbg_0_n_39_15));
  XNOR2_X1_LVT dbg_0_i_39_32 (.ZN(dbg_0_n_71), .A(dbg_0_mem_cnt[15]), .B(
      dbg_0_n_39_16));
  AOI22_X1_LVT dbg_0_i_40_31 (.ZN(dbg_0_n_40_16), .A1(dbg_0_n_40_0), .A2(
      dbg_0_n_71), .B1(dbg_0_n_102), .B2(dbg_0_dbg_din[15]));
  INV_X1_LVT dbg_0_i_40_32 (.ZN(dbg_0_n_87), .A(dbg_0_n_40_16));
  DFFR_X1_LVT \dbg_0_mem_cnt_reg[15] (.Q(dbg_0_mem_cnt[15]), .QN(), .CK(dbg_clk), 
      .D(dbg_0_n_87), .RN(dbg_0_n_104));
  NOR4_X1_LVT dbg_0_i_37_3 (.ZN(dbg_0_n_37_3), .A1(dbg_0_mem_cnt[12]), .A2(
      dbg_0_mem_cnt[13]), .A3(dbg_0_mem_cnt[14]), .A4(dbg_0_mem_cnt[15]));
  NAND4_X1_LVT dbg_0_i_37_4 (.ZN(dbg_0_n_37_4), .A1(dbg_0_n_37_0), .A2(
      dbg_0_n_37_1), .A3(dbg_0_n_37_2), .A4(dbg_0_n_37_3));
  CLKGATETST_X1_LVT dbg_0_clk_gate_mem_ctl_reg (.GCK(dbg_0_n_2), .CK(dbg_clk), 
      .E(dbg_0_mem_ctl_wr), .SE(1'b0));
  DFFR_X1_LVT \dbg_0_mem_ctl_reg[1] (.Q(dbg_0_mem_ctl[0]), .QN(), .CK(dbg_0_n_2), 
      .D(dbg_0_dbg_din[1]), .RN(dbg_0_n_104));
  OAI21_X1_LVT dbg_0_i_6_0 (.ZN(dbg_0_n_6_0), .A(dbg_0_mem_burst), .B1(
      dbg_0_dbg_wr), .B2(dbg_0_dbg_rd));
  INV_X1_LVT dbg_0_i_4_0 (.ZN(dbg_0_n_3), .A(dbg_0_mem_ctl[0]));
  AND2_X1_LVT dbg_0_i_5_0 (.ZN(dbg_0_mem_burst_rd), .A1(dbg_0_n_3), .A2(
      dbg_0_mem_burst_start));
  INV_X1_LVT dbg_0_i_6_1 (.ZN(dbg_0_n_6_1), .A(dbg_0_mem_burst_rd));
  NAND2_X1_LVT dbg_0_i_6_2 (.ZN(dbg_0_n_4), .A1(dbg_0_n_6_0), .A2(dbg_0_n_6_1));
  DFFR_X1_LVT dbg_0_mem_startb_reg (.Q(dbg_0_mem_startb), .QN(), .CK(dbg_clk), 
      .D(dbg_0_n_4), .RN(dbg_0_n_104));
  NOR4_X1_LVT dbg_0_i_0_0 (.ZN(dbg_0_n_0_0), .A1(dbg_0_mem_cnt[0]), .A2(
      dbg_0_mem_cnt[1]), .A3(dbg_0_mem_cnt[2]), .A4(dbg_0_mem_cnt[3]));
  NOR4_X1_LVT dbg_0_i_0_1 (.ZN(dbg_0_n_0_1), .A1(dbg_0_mem_cnt[4]), .A2(
      dbg_0_mem_cnt[5]), .A3(dbg_0_mem_cnt[6]), .A4(dbg_0_mem_cnt[7]));
  NOR4_X1_LVT dbg_0_i_0_2 (.ZN(dbg_0_n_0_2), .A1(dbg_0_mem_cnt[8]), .A2(
      dbg_0_mem_cnt[9]), .A3(dbg_0_mem_cnt[10]), .A4(dbg_0_mem_cnt[11]));
  NOR4_X1_LVT dbg_0_i_0_3 (.ZN(dbg_0_n_0_3), .A1(dbg_0_mem_cnt[12]), .A2(
      dbg_0_mem_cnt[13]), .A3(dbg_0_mem_cnt[14]), .A4(dbg_0_mem_cnt[15]));
  AND4_X1_LVT dbg_0_i_0_4 (.ZN(dbg_0_n_0), .A1(dbg_0_n_0_0), .A2(dbg_0_n_0_1), 
      .A3(dbg_0_n_0_2), .A4(dbg_0_n_0_3));
  AOI21_X1_LVT dbg_0_i_8_0 (.ZN(dbg_0_n_8_0), .A(dbg_0_mem_startb), .B1(
      dbg_0_n_0), .B2(dbg_0_mem_start));
  INV_X1_LVT dbg_0_i_8_1 (.ZN(dbg_0_n_5), .A(dbg_0_n_8_0));
  NAND2_X1_LVT dbg_0_i_9_0 (.ZN(dbg_0_n_9_0), .A1(cpu_halt_st), .A2(dbg_0_n_5));
  INV_X1_LVT dbg_0_i_9_1 (.ZN(dbg_0_n_9_1), .A(dbg_0_n_9_0));
  INV_X1_LVT dbg_0_i_9_7 (.ZN(dbg_0_n_9_6), .A(cpu_halt_st));
  AOI21_X1_LVT dbg_0_i_9_2 (.ZN(dbg_0_n_9_2), .A(dbg_0_n_9_1), .B1(dbg_0_n_9_6), 
      .B2(dbg_0_n_5));
  INV_X1_LVT dbg_0_i_9_4 (.ZN(dbg_0_n_9_4), .A(dbg_0_mem_state[1]));
  NAND2_X1_LVT dbg_0_i_9_5 (.ZN(dbg_0_n_9_5), .A1(dbg_0_n_9_4), .A2(
      dbg_0_mem_state[0]));
  OAI22_X1_LVT dbg_0_i_9_8 (.ZN(dbg_0_mem_state_nxt_reg[1]), .A1(dbg_0_n_9_3), 
      .A2(dbg_0_n_9_0), .B1(dbg_0_n_9_5), .B2(dbg_0_n_9_6));
  DFFR_X1_LVT \dbg_0_mem_state_reg[1] (.Q(dbg_0_mem_state[1]), .QN(), .CK(
      dbg_clk), .D(dbg_0_mem_state_nxt_reg[1]), .RN(dbg_0_n_104));
  OR2_X1_LVT dbg_0_i_9_3 (.ZN(dbg_0_n_9_3), .A1(dbg_0_mem_state[0]), .A2(
      dbg_0_mem_state[1]));
  OAI22_X1_LVT dbg_0_i_9_6 (.ZN(dbg_0_mem_state_nxt_reg[0]), .A1(dbg_0_n_9_2), 
      .A2(dbg_0_n_9_3), .B1(dbg_0_n_9_5), .B2(cpu_halt_st));
  DFFR_X1_LVT \dbg_0_mem_state_reg[0] (.Q(dbg_0_mem_state[0]), .QN(), .CK(dbg_clk), 
      .D(dbg_0_mem_state_nxt_reg[0]), .RN(dbg_0_n_104));
  AND2_X1_LVT dbg_0_i_12_0 (.ZN(dbg_0_n_6), .A1(dbg_0_mem_state[0]), .A2(
      dbg_0_mem_state[1]));
  INV_X1_LVT dbg_0_i_12_1 (.ZN(dbg_0_n_12_0), .A(dbg_0_mem_state[1]));
  NOR2_X1_LVT dbg_0_i_12_2 (.ZN(dbg_0_n_7), .A1(dbg_0_n_12_0), .A2(
      dbg_0_mem_state[0]));
  OR2_X1_LVT dbg_0_i_13_0 (.ZN(dbg_0_mem_access), .A1(dbg_0_n_6), .A2(dbg_0_n_7));
  DFFR_X1_LVT \dbg_0_mem_ctl_reg[2] (.Q(dbg_0_mem_ctl[1]), .QN(), .CK(dbg_0_n_2), 
      .D(dbg_0_dbg_din[2]), .RN(dbg_0_n_104));
  INV_X1_LVT dbg_0_i_23_0 (.ZN(dbg_0_n_47), .A(dbg_0_mem_ctl[1]));
  AND2_X1_LVT dbg_0_i_24_0 (.ZN(dbg_mem_en), .A1(dbg_0_mem_access), .A2(
      dbg_0_n_47));
  AND2_X1_LVT dbg_0_i_25_0 (.ZN(dbg_0_n_48), .A1(dbg_0_mem_ctl[0]), .A2(
      dbg_mem_en));
  NOR2_X1_LVT dbg_0_i_49_3 (.ZN(dbg_0_n_49_3), .A1(dbg_0_n_49_0), .A2(
      dbg_0_dbg_addr_in[1]));
  NAND2_X1_LVT dbg_0_i_49_12 (.ZN(dbg_0_n_49_12), .A1(dbg_0_n_49_3), .A2(
      dbg_0_dbg_addr_in[2]));
  NOR2_X1_LVT dbg_0_i_49_27 (.ZN(dbg_0_n_96), .A1(dbg_0_n_49_12), .A2(
      dbg_0_n_49_20));
  AND2_X1_LVT dbg_0_i_50_3 (.ZN(dbg_0_n_101), .A1(dbg_0_dbg_wr), .A2(dbg_0_n_96));
  INV_X1_LVT dbg_0_i_20_0 (.ZN(dbg_0_n_20_0), .A(dbg_0_n_101));
  NOR4_X1_LVT dbg_0_i_17_0 (.ZN(dbg_0_n_17_0), .A1(dbg_0_mem_cnt[0]), .A2(
      dbg_0_mem_cnt[1]), .A3(dbg_0_mem_cnt[2]), .A4(dbg_0_mem_cnt[3]));
  NOR4_X1_LVT dbg_0_i_17_1 (.ZN(dbg_0_n_17_1), .A1(dbg_0_mem_cnt[4]), .A2(
      dbg_0_mem_cnt[5]), .A3(dbg_0_mem_cnt[6]), .A4(dbg_0_mem_cnt[7]));
  NOR4_X1_LVT dbg_0_i_17_2 (.ZN(dbg_0_n_17_2), .A1(dbg_0_mem_cnt[8]), .A2(
      dbg_0_mem_cnt[9]), .A3(dbg_0_mem_cnt[10]), .A4(dbg_0_mem_cnt[11]));
  NOR4_X1_LVT dbg_0_i_17_3 (.ZN(dbg_0_n_17_3), .A1(dbg_0_mem_cnt[12]), .A2(
      dbg_0_mem_cnt[13]), .A3(dbg_0_mem_cnt[14]), .A4(dbg_0_mem_cnt[15]));
  NAND4_X1_LVT dbg_0_i_17_4 (.ZN(dbg_0_n_17_4), .A1(dbg_0_n_17_0), .A2(
      dbg_0_n_17_1), .A3(dbg_0_n_17_2), .A4(dbg_0_n_17_3));
  INV_X1_LVT dbg_0_i_16_0 (.ZN(dbg_0_n_16_0), .A(dbg_0_dbg_mem_acc));
  DFFR_X1_LVT \dbg_0_mem_ctl_reg[3] (.Q(dbg_0_mem_ctl[2]), .QN(), .CK(dbg_0_n_2), 
      .D(dbg_0_dbg_din[3]), .RN(dbg_0_n_104));
  NOR2_X1_LVT dbg_0_i_16_1 (.ZN(dbg_0_n_10), .A1(dbg_0_n_16_0), .A2(
      dbg_0_mem_ctl[2]));
  NAND2_X1_LVT dbg_0_i_17_5 (.ZN(dbg_0_n_17_5), .A1(dbg_0_n_10), .A2(
      dbg_0_mem_burst));
  AND4_X1_LVT dbg_0_i_17_6 (.ZN(dbg_0_n_11), .A1(dbg_0_n_17_4), .A2(dbg_0_n_17_5), 
      .A3(dbg_0_mem_burst), .A4(dbg_0_n_53));
  HA_X1_LVT dbg_0_i_19_0 (.CO(dbg_0_n_19_0), .S(dbg_0_n_13), .A(dbg_0_n_11), .B(
      dbg_mem_addr[0]));
  AOI22_X1_LVT dbg_0_i_20_1 (.ZN(dbg_0_n_20_1), .A1(dbg_0_n_20_0), .A2(
      dbg_0_n_13), .B1(dbg_0_dbg_din[0]), .B2(dbg_0_n_101));
  INV_X1_LVT dbg_0_i_20_2 (.ZN(dbg_0_n_29), .A(dbg_0_n_20_1));
  DFFR_X1_LVT \dbg_0_mem_addr_reg[0] (.Q(dbg_mem_addr[0]), .QN(), .CK(dbg_clk), 
      .D(dbg_0_n_29), .RN(dbg_0_n_104));
  NAND2_X1_LVT dbg_0_i_22_2 (.ZN(dbg_0_n_46), .A1(dbg_mem_addr[0]), .A2(
      dbg_0_mem_ctl[2]));
  AND2_X1_LVT dbg_0_i_26_0 (.ZN(dbg_mem_wr[0]), .A1(dbg_0_n_48), .A2(dbg_0_n_46));
  INV_X1_LVT dbg_0_i_22_0 (.ZN(dbg_0_n_22_0), .A(dbg_mem_addr[0]));
  NAND2_X1_LVT dbg_0_i_22_1 (.ZN(dbg_0_n_45), .A1(dbg_0_n_22_0), .A2(
      dbg_0_mem_ctl[2]));
  AND2_X1_LVT dbg_0_i_26_1 (.ZN(dbg_mem_wr[1]), .A1(dbg_0_n_48), .A2(dbg_0_n_45));
  OR2_X1_LVT dbg_0_i_27_0 (.ZN(dbg_0_n_49), .A1(dbg_mem_wr[0]), .A2(dbg_mem_wr[1]));
  OR2_X1_LVT dbg_0_i_31_0 (.ZN(dbg_0_n_51), .A1(dbg_0_mem_burst), .A2(
      dbg_0_mem_burst_rd));
  INV_X1_LVT dbg_0_i_32_0 (.ZN(dbg_0_n_32_0), .A(dbg_0_n_51));
  AND2_X1_LVT dbg_0_i_14_0 (.ZN(dbg_0_n_9), .A1(dbg_0_mem_ctl[1]), .A2(
      dbg_0_mem_access));
  AND2_X1_LVT dbg_0_i_28_0 (.ZN(dbg_0_dbg_reg_rd), .A1(dbg_0_n_3), .A2(dbg_0_n_9));
  AND2_X1_LVT dbg_0_i_29_0 (.ZN(dbg_0_dbg_mem_rd), .A1(dbg_0_n_3), .A2(
      dbg_mem_en));
  DFFR_X1_LVT dbg_0_dbg_mem_rd_dly_reg (.Q(dbg_0_dbg_mem_rd_dly), .QN(), .CK(
      dbg_clk), .D(dbg_0_dbg_mem_rd), .RN(dbg_0_n_104));
  OR2_X1_LVT dbg_0_i_30_0 (.ZN(dbg_0_n_50), .A1(dbg_0_dbg_reg_rd), .A2(
      dbg_0_dbg_mem_rd_dly));
  AOI22_X1_LVT dbg_0_i_32_1 (.ZN(dbg_0_n_32_1), .A1(dbg_0_n_32_0), .A2(
      dbg_0_dbg_rd), .B1(dbg_0_n_50), .B2(dbg_0_n_51));
  INV_X1_LVT dbg_0_i_32_2 (.ZN(dbg_0_n_52), .A(dbg_0_n_32_1));
  DFFR_X1_LVT dbg_0_dbg_rd_rdy_reg (.Q(dbg_0_dbg_rd_rdy), .QN(), .CK(dbg_clk), 
      .D(dbg_0_n_52), .RN(dbg_0_n_104));
  AOI21_X1_LVT dbg_0_i_34_0 (.ZN(dbg_0_n_34_0), .A(dbg_0_n_49), .B1(
      dbg_0_dbg_rd_rdy), .B2(dbg_0_n_47));
  INV_X1_LVT dbg_0_i_34_1 (.ZN(dbg_0_dbg_mem_acc), .A(dbg_0_n_34_0));
  AND2_X1_LVT dbg_0_i_15_0 (.ZN(dbg_reg_wr), .A1(dbg_0_mem_ctl[0]), .A2(dbg_0_n_9));
  NOR2_X1_LVT dbg_0_i_35_0 (.ZN(dbg_0_n_35_0), .A1(dbg_0_dbg_mem_acc), .A2(
      dbg_reg_wr));
  NAND2_X1_LVT dbg_0_i_35_1 (.ZN(dbg_0_n_35_1), .A1(dbg_0_mem_ctl[1]), .A2(
      dbg_0_dbg_rd_rdy));
  NAND2_X1_LVT dbg_0_i_35_2 (.ZN(dbg_0_n_53), .A1(dbg_0_n_35_0), .A2(
      dbg_0_n_35_1));
  AND2_X1_LVT dbg_0_i_36_0 (.ZN(dbg_0_n_54), .A1(dbg_0_n_53), .A2(
      dbg_0_mem_burst));
  AND2_X1_LVT dbg_0_i_37_5 (.ZN(dbg_0_n_55), .A1(dbg_0_n_37_4), .A2(dbg_0_n_54));
  XNOR2_X1_LVT dbg_0_i_39_0 (.ZN(dbg_0_n_39_0), .A(dbg_0_n_55), .B(
      dbg_0_mem_cnt[0]));
  INV_X1_LVT dbg_0_i_39_1 (.ZN(dbg_0_n_56), .A(dbg_0_n_39_0));
  AOI22_X1_LVT dbg_0_i_40_1 (.ZN(dbg_0_n_40_1), .A1(dbg_0_n_40_0), .A2(
      dbg_0_n_56), .B1(dbg_0_dbg_din[0]), .B2(dbg_0_n_102));
  INV_X1_LVT dbg_0_i_40_2 (.ZN(dbg_0_n_72), .A(dbg_0_n_40_1));
  DFFR_X1_LVT \dbg_0_mem_cnt_reg[0] (.Q(dbg_0_mem_cnt[0]), .QN(), .CK(dbg_clk), 
      .D(dbg_0_n_72), .RN(dbg_0_n_104));
  NOR4_X1_LVT dbg_0_i_42_0 (.ZN(dbg_0_n_42_0), .A1(dbg_0_mem_cnt[0]), .A2(
      dbg_0_mem_cnt[1]), .A3(dbg_0_mem_cnt[2]), .A4(dbg_0_mem_cnt[3]));
  NOR4_X1_LVT dbg_0_i_42_1 (.ZN(dbg_0_n_42_1), .A1(dbg_0_mem_cnt[4]), .A2(
      dbg_0_mem_cnt[5]), .A3(dbg_0_mem_cnt[6]), .A4(dbg_0_mem_cnt[7]));
  NOR4_X1_LVT dbg_0_i_42_2 (.ZN(dbg_0_n_42_2), .A1(dbg_0_mem_cnt[8]), .A2(
      dbg_0_mem_cnt[9]), .A3(dbg_0_mem_cnt[10]), .A4(dbg_0_mem_cnt[11]));
  NOR4_X1_LVT dbg_0_i_42_3 (.ZN(dbg_0_n_42_3), .A1(dbg_0_mem_cnt[12]), .A2(
      dbg_0_mem_cnt[13]), .A3(dbg_0_mem_cnt[14]), .A4(dbg_0_mem_cnt[15]));
  NAND4_X1_LVT dbg_0_i_42_4 (.ZN(dbg_0_n_88), .A1(dbg_0_n_42_0), .A2(
      dbg_0_n_42_1), .A3(dbg_0_n_42_2), .A4(dbg_0_n_42_3));
  AND2_X1_LVT dbg_0_i_43_0 (.ZN(dbg_0_mem_burst_start), .A1(dbg_0_mem_start), 
      .A2(dbg_0_n_88));
  OAI21_X1_LVT dbg_0_i_44_0 (.ZN(dbg_0_n_44_0), .A(dbg_0_n_0), .B1(dbg_0_dbg_wr), 
      .B2(dbg_0_dbg_rd_rdy));
  INV_X1_LVT dbg_0_i_44_1 (.ZN(dbg_0_mem_burst_end), .A(dbg_0_n_44_0));
  INV_X1_LVT dbg_0_i_46_1 (.ZN(dbg_0_n_46_1), .A(dbg_0_mem_burst_end));
  INV_X1_LVT dbg_0_i_46_0 (.ZN(dbg_0_n_46_0), .A(dbg_0_mem_burst_start));
  NAND2_X1_LVT dbg_0_i_46_2 (.ZN(dbg_0_n_90), .A1(dbg_0_n_46_1), .A2(
      dbg_0_n_46_0));
  CLKGATETST_X1_LVT dbg_0_clk_gate_mem_burst_reg (.GCK(dbg_0_n_89), .CK(dbg_clk), 
      .E(dbg_0_n_90), .SE(1'b0));
  DFFR_X1_LVT dbg_0_mem_burst_reg (.Q(dbg_0_mem_burst), .QN(), .CK(dbg_0_n_89), 
      .D(dbg_0_mem_burst_start), .RN(dbg_0_n_104));
  INV_X1_LVT dbg_0_i_48_0 (.ZN(dbg_0_n_48_0), .A(dbg_0_mem_burst));
  AND2_X1_LVT dbg_0_i_48_1 (.ZN(dbg_0_dbg_addr_in[0]), .A1(dbg_0_n_48_0), .A2(
      dbg_0_dbg_addr[0]));
  INV_X1_LVT dbg_0_i_49_0 (.ZN(dbg_0_n_49_0), .A(dbg_0_dbg_addr_in[0]));
  INV_X1_LVT dbg_0_i_49_1 (.ZN(dbg_0_n_49_1), .A(dbg_0_dbg_addr_in[1]));
  NOR2_X1_LVT dbg_0_i_49_5 (.ZN(dbg_0_n_49_5), .A1(dbg_0_n_49_0), .A2(
      dbg_0_n_49_1));
  NAND2_X1_LVT dbg_0_i_49_14 (.ZN(dbg_0_n_49_14), .A1(dbg_0_n_49_5), .A2(
      dbg_0_dbg_addr_in[2]));
  NOR2_X1_LVT dbg_0_i_49_29 (.ZN(dbg_0_n_98), .A1(dbg_0_n_49_14), .A2(
      dbg_0_n_49_20));
  NAND2_X1_LVT dbg_0_i_78_125 (.ZN(dbg_0_n_78_110), .A1(dbg_0_n_98), .A2(
      dbg_0_mem_cnt[15]));
  AOI22_X1_LVT dbg_0_i_20_29 (.ZN(dbg_0_n_20_15), .A1(dbg_0_n_20_0), .A2(
      dbg_0_n_27), .B1(dbg_0_n_101), .B2(dbg_0_dbg_din[14]));
  INV_X1_LVT dbg_0_i_20_30 (.ZN(dbg_0_n_43), .A(dbg_0_n_20_15));
  DFFR_X1_LVT \dbg_0_mem_addr_reg[14] (.Q(dbg_mem_addr[14]), .QN(), .CK(dbg_clk), 
      .D(dbg_0_n_43), .RN(dbg_0_n_104));
  AOI22_X1_LVT dbg_0_i_20_27 (.ZN(dbg_0_n_20_14), .A1(dbg_0_n_20_0), .A2(
      dbg_0_n_26), .B1(dbg_0_n_101), .B2(dbg_0_dbg_din[13]));
  INV_X1_LVT dbg_0_i_20_28 (.ZN(dbg_0_n_42), .A(dbg_0_n_20_14));
  DFFR_X1_LVT \dbg_0_mem_addr_reg[13] (.Q(dbg_mem_addr[13]), .QN(), .CK(dbg_clk), 
      .D(dbg_0_n_42), .RN(dbg_0_n_104));
  AOI22_X1_LVT dbg_0_i_20_25 (.ZN(dbg_0_n_20_13), .A1(dbg_0_n_20_0), .A2(
      dbg_0_n_25), .B1(dbg_0_n_101), .B2(dbg_0_dbg_din[12]));
  INV_X1_LVT dbg_0_i_20_26 (.ZN(dbg_0_n_41), .A(dbg_0_n_20_13));
  DFFR_X1_LVT \dbg_0_mem_addr_reg[12] (.Q(dbg_mem_addr[12]), .QN(), .CK(dbg_clk), 
      .D(dbg_0_n_41), .RN(dbg_0_n_104));
  AOI22_X1_LVT dbg_0_i_20_23 (.ZN(dbg_0_n_20_12), .A1(dbg_0_n_20_0), .A2(
      dbg_0_n_24), .B1(dbg_0_n_101), .B2(dbg_0_dbg_din[11]));
  INV_X1_LVT dbg_0_i_20_24 (.ZN(dbg_0_n_40), .A(dbg_0_n_20_12));
  DFFR_X1_LVT \dbg_0_mem_addr_reg[11] (.Q(dbg_mem_addr[11]), .QN(), .CK(dbg_clk), 
      .D(dbg_0_n_40), .RN(dbg_0_n_104));
  AOI22_X1_LVT dbg_0_i_20_21 (.ZN(dbg_0_n_20_11), .A1(dbg_0_n_20_0), .A2(
      dbg_0_n_23), .B1(dbg_0_n_101), .B2(dbg_0_dbg_din[10]));
  INV_X1_LVT dbg_0_i_20_22 (.ZN(dbg_0_n_39), .A(dbg_0_n_20_11));
  DFFR_X1_LVT \dbg_0_mem_addr_reg[10] (.Q(dbg_mem_addr[10]), .QN(), .CK(dbg_clk), 
      .D(dbg_0_n_39), .RN(dbg_0_n_104));
  AOI22_X1_LVT dbg_0_i_20_19 (.ZN(dbg_0_n_20_10), .A1(dbg_0_n_20_0), .A2(
      dbg_0_n_22), .B1(dbg_0_n_101), .B2(dbg_0_dbg_din[9]));
  INV_X1_LVT dbg_0_i_20_20 (.ZN(dbg_0_n_38), .A(dbg_0_n_20_10));
  DFFR_X1_LVT \dbg_0_mem_addr_reg[9] (.Q(dbg_mem_addr[9]), .QN(), .CK(dbg_clk), 
      .D(dbg_0_n_38), .RN(dbg_0_n_104));
  AOI22_X1_LVT dbg_0_i_20_17 (.ZN(dbg_0_n_20_9), .A1(dbg_0_n_20_0), .A2(
      dbg_0_n_21), .B1(dbg_0_n_101), .B2(dbg_0_dbg_din[8]));
  INV_X1_LVT dbg_0_i_20_18 (.ZN(dbg_0_n_37), .A(dbg_0_n_20_9));
  DFFR_X1_LVT \dbg_0_mem_addr_reg[8] (.Q(dbg_mem_addr[8]), .QN(), .CK(dbg_clk), 
      .D(dbg_0_n_37), .RN(dbg_0_n_104));
  AOI22_X1_LVT dbg_0_i_20_15 (.ZN(dbg_0_n_20_8), .A1(dbg_0_n_20_0), .A2(
      dbg_0_n_20), .B1(dbg_0_n_101), .B2(dbg_0_dbg_din[7]));
  INV_X1_LVT dbg_0_i_20_16 (.ZN(dbg_0_n_36), .A(dbg_0_n_20_8));
  DFFR_X1_LVT \dbg_0_mem_addr_reg[7] (.Q(dbg_mem_addr[7]), .QN(), .CK(dbg_clk), 
      .D(dbg_0_n_36), .RN(dbg_0_n_104));
  AOI22_X1_LVT dbg_0_i_20_13 (.ZN(dbg_0_n_20_7), .A1(dbg_0_n_20_0), .A2(
      dbg_0_n_19), .B1(dbg_0_n_101), .B2(dbg_0_dbg_din[6]));
  INV_X1_LVT dbg_0_i_20_14 (.ZN(dbg_0_n_35), .A(dbg_0_n_20_7));
  DFFR_X1_LVT \dbg_0_mem_addr_reg[6] (.Q(dbg_mem_addr[6]), .QN(), .CK(dbg_clk), 
      .D(dbg_0_n_35), .RN(dbg_0_n_104));
  AOI22_X1_LVT dbg_0_i_20_11 (.ZN(dbg_0_n_20_6), .A1(dbg_0_n_20_0), .A2(
      dbg_0_n_18), .B1(dbg_0_n_101), .B2(dbg_0_dbg_din[5]));
  INV_X1_LVT dbg_0_i_20_12 (.ZN(dbg_0_n_34), .A(dbg_0_n_20_6));
  DFFR_X1_LVT \dbg_0_mem_addr_reg[5] (.Q(dbg_mem_addr[5]), .QN(), .CK(dbg_clk), 
      .D(dbg_0_n_34), .RN(dbg_0_n_104));
  AOI22_X1_LVT dbg_0_i_20_9 (.ZN(dbg_0_n_20_5), .A1(dbg_0_n_20_0), .A2(
      dbg_0_n_17), .B1(dbg_0_n_101), .B2(dbg_0_dbg_din[4]));
  INV_X1_LVT dbg_0_i_20_10 (.ZN(dbg_0_n_33), .A(dbg_0_n_20_5));
  DFFR_X1_LVT \dbg_0_mem_addr_reg[4] (.Q(dbg_mem_addr[4]), .QN(), .CK(dbg_clk), 
      .D(dbg_0_n_33), .RN(dbg_0_n_104));
  AOI22_X1_LVT dbg_0_i_20_7 (.ZN(dbg_0_n_20_4), .A1(dbg_0_n_20_0), .A2(
      dbg_0_n_16), .B1(dbg_0_n_101), .B2(dbg_0_dbg_din[3]));
  INV_X1_LVT dbg_0_i_20_8 (.ZN(dbg_0_n_32), .A(dbg_0_n_20_4));
  DFFR_X1_LVT \dbg_0_mem_addr_reg[3] (.Q(dbg_mem_addr[3]), .QN(), .CK(dbg_clk), 
      .D(dbg_0_n_32), .RN(dbg_0_n_104));
  AOI22_X1_LVT dbg_0_i_20_5 (.ZN(dbg_0_n_20_3), .A1(dbg_0_n_20_0), .A2(
      dbg_0_n_15), .B1(dbg_0_n_101), .B2(dbg_0_dbg_din[2]));
  INV_X1_LVT dbg_0_i_20_6 (.ZN(dbg_0_n_31), .A(dbg_0_n_20_3));
  DFFR_X1_LVT \dbg_0_mem_addr_reg[2] (.Q(dbg_mem_addr[2]), .QN(), .CK(dbg_clk), 
      .D(dbg_0_n_31), .RN(dbg_0_n_104));
  INV_X1_LVT dbg_0_i_17_7 (.ZN(dbg_0_n_17_6), .A(dbg_0_n_17_4));
  NOR2_X1_LVT dbg_0_i_17_8 (.ZN(dbg_0_n_12), .A1(dbg_0_n_17_6), .A2(dbg_0_n_17_5));
  AOI22_X1_LVT dbg_0_i_20_3 (.ZN(dbg_0_n_20_2), .A1(dbg_0_n_20_0), .A2(
      dbg_0_n_14), .B1(dbg_0_n_101), .B2(dbg_0_dbg_din[1]));
  INV_X1_LVT dbg_0_i_20_4 (.ZN(dbg_0_n_30), .A(dbg_0_n_20_2));
  DFFR_X1_LVT \dbg_0_mem_addr_reg[1] (.Q(dbg_mem_addr[1]), .QN(), .CK(dbg_clk), 
      .D(dbg_0_n_30), .RN(dbg_0_n_104));
  FA_X1_LVT dbg_0_i_19_1 (.CO(dbg_0_n_19_1), .S(dbg_0_n_14), .A(dbg_0_n_12), .B(
      dbg_mem_addr[1]), .CI(dbg_0_n_19_0));
  HA_X1_LVT dbg_0_i_19_2 (.CO(dbg_0_n_19_2), .S(dbg_0_n_15), .A(dbg_mem_addr[2]), 
      .B(dbg_0_n_19_1));
  HA_X1_LVT dbg_0_i_19_3 (.CO(dbg_0_n_19_3), .S(dbg_0_n_16), .A(dbg_mem_addr[3]), 
      .B(dbg_0_n_19_2));
  HA_X1_LVT dbg_0_i_19_4 (.CO(dbg_0_n_19_4), .S(dbg_0_n_17), .A(dbg_mem_addr[4]), 
      .B(dbg_0_n_19_3));
  HA_X1_LVT dbg_0_i_19_5 (.CO(dbg_0_n_19_5), .S(dbg_0_n_18), .A(dbg_mem_addr[5]), 
      .B(dbg_0_n_19_4));
  HA_X1_LVT dbg_0_i_19_6 (.CO(dbg_0_n_19_6), .S(dbg_0_n_19), .A(dbg_mem_addr[6]), 
      .B(dbg_0_n_19_5));
  HA_X1_LVT dbg_0_i_19_7 (.CO(dbg_0_n_19_7), .S(dbg_0_n_20), .A(dbg_mem_addr[7]), 
      .B(dbg_0_n_19_6));
  HA_X1_LVT dbg_0_i_19_8 (.CO(dbg_0_n_19_8), .S(dbg_0_n_21), .A(dbg_mem_addr[8]), 
      .B(dbg_0_n_19_7));
  HA_X1_LVT dbg_0_i_19_9 (.CO(dbg_0_n_19_9), .S(dbg_0_n_22), .A(dbg_mem_addr[9]), 
      .B(dbg_0_n_19_8));
  HA_X1_LVT dbg_0_i_19_10 (.CO(dbg_0_n_19_10), .S(dbg_0_n_23), .A(
      dbg_mem_addr[10]), .B(dbg_0_n_19_9));
  HA_X1_LVT dbg_0_i_19_11 (.CO(dbg_0_n_19_11), .S(dbg_0_n_24), .A(
      dbg_mem_addr[11]), .B(dbg_0_n_19_10));
  HA_X1_LVT dbg_0_i_19_12 (.CO(dbg_0_n_19_12), .S(dbg_0_n_25), .A(
      dbg_mem_addr[12]), .B(dbg_0_n_19_11));
  HA_X1_LVT dbg_0_i_19_13 (.CO(dbg_0_n_19_13), .S(dbg_0_n_26), .A(
      dbg_mem_addr[13]), .B(dbg_0_n_19_12));
  HA_X1_LVT dbg_0_i_19_14 (.CO(dbg_0_n_19_14), .S(dbg_0_n_27), .A(
      dbg_mem_addr[14]), .B(dbg_0_n_19_13));
  XNOR2_X1_LVT dbg_0_i_19_15 (.ZN(dbg_0_n_19_15), .A(dbg_mem_addr[15]), .B(
      dbg_0_n_19_14));
  INV_X1_LVT dbg_0_i_19_16 (.ZN(dbg_0_n_28), .A(dbg_0_n_19_15));
  AOI22_X1_LVT dbg_0_i_20_31 (.ZN(dbg_0_n_20_16), .A1(dbg_0_n_20_0), .A2(
      dbg_0_n_28), .B1(dbg_0_n_101), .B2(dbg_0_dbg_din[15]));
  INV_X1_LVT dbg_0_i_20_32 (.ZN(dbg_0_n_44), .A(dbg_0_n_20_16));
  DFFR_X1_LVT \dbg_0_mem_addr_reg[15] (.Q(dbg_mem_addr[15]), .QN(), .CK(dbg_clk), 
      .D(dbg_0_n_44), .RN(dbg_0_n_104));
  NAND2_X1_LVT dbg_0_i_78_126 (.ZN(dbg_0_n_78_111), .A1(dbg_0_n_96), .A2(
      dbg_mem_addr[15]));
  NOR2_X1_LVT dbg_0_i_49_4 (.ZN(dbg_0_n_49_4), .A1(dbg_0_dbg_addr_in[0]), .A2(
      dbg_0_n_49_1));
  NAND2_X1_LVT dbg_0_i_49_13 (.ZN(dbg_0_n_49_13), .A1(dbg_0_n_49_4), .A2(
      dbg_0_dbg_addr_in[2]));
  NOR2_X1_LVT dbg_0_i_49_28 (.ZN(dbg_0_n_97), .A1(dbg_0_n_49_13), .A2(
      dbg_0_n_49_20));
  AND2_X1_LVT dbg_0_i_50_4 (.ZN(dbg_0_mem_data_wr), .A1(dbg_0_dbg_wr), .A2(
      dbg_0_n_97));
  INV_X1_LVT dbg_0_i_70_1 (.ZN(dbg_0_n_70_0), .A(dbg_0_dbg_reg_rd));
  NOR2_X1_LVT dbg_0_i_70_2 (.ZN(dbg_0_n_136), .A1(dbg_0_n_70_0), .A2(
      dbg_0_mem_data_wr));
  NOR2_X1_LVT dbg_0_i_70_0 (.ZN(dbg_0_n_135), .A1(dbg_0_dbg_reg_rd), .A2(
      dbg_0_mem_data_wr));
  INV_X1_LVT dbg_0_i_67_0 (.ZN(dbg_0_n_115), .A(dbg_0_mem_ctl[2]));
  AND2_X1_LVT dbg_0_i_68_24 (.ZN(dbg_0_n_133), .A1(dbg_0_n_115), .A2(
      dbg_mem_din[15]));
  AOI222_X1_LVT dbg_0_i_71_30 (.ZN(dbg_0_n_71_15), .A1(dbg_0_mem_data_wr), .A2(
      dbg_0_dbg_din[15]), .B1(dbg_0_n_136), .B2(dbg_reg_din[15]), .C1(
      dbg_0_n_135), .C2(dbg_0_n_133));
  INV_X1_LVT dbg_0_i_71_31 (.ZN(dbg_0_n_152), .A(dbg_0_n_71_15));
  INV_X1_LVT dbg_0_i_72_0 (.ZN(dbg_0_n_72_0), .A(dbg_0_dbg_reg_rd));
  INV_X1_LVT dbg_0_i_72_1 (.ZN(dbg_0_n_72_1), .A(dbg_0_mem_data_wr));
  NAND3_X1_LVT dbg_0_i_72_2 (.ZN(dbg_0_n_72_2), .A1(dbg_0_n_72_0), .A2(
      dbg_0_n_72_1), .A3(dbg_0_dbg_mem_rd_dly));
  NAND3_X1_LVT dbg_0_i_72_3 (.ZN(dbg_0_n_153), .A1(dbg_0_n_72_2), .A2(
      dbg_0_n_72_0), .A3(dbg_0_n_72_1));
  CLKGATETST_X1_LVT dbg_0_clk_gate_mem_data_reg (.GCK(dbg_0_n_134), .CK(dbg_clk), 
      .E(dbg_0_n_153), .SE(1'b0));
  DFFR_X1_LVT \dbg_0_mem_data_reg[15] (.Q(dbg_0_mem_data[15]), .QN(), .CK(
      dbg_0_n_134), .D(dbg_0_n_152), .RN(dbg_0_n_104));
  NAND2_X1_LVT dbg_0_i_78_127 (.ZN(dbg_0_n_78_112), .A1(dbg_0_n_97), .A2(
      dbg_0_mem_data[15]));
  INV_X1_LVT dbg_0_i_49_6 (.ZN(dbg_0_n_49_6), .A(dbg_0_dbg_addr_in[2]));
  NAND2_X1_LVT dbg_0_i_49_8 (.ZN(dbg_0_n_49_8), .A1(dbg_0_n_49_3), .A2(
      dbg_0_n_49_6));
  NOR2_X1_LVT dbg_0_i_49_23 (.ZN(dbg_0_n_92), .A1(dbg_0_n_49_8), .A2(
      dbg_0_n_49_20));
  NAND2_X1_LVT dbg_0_i_78_128 (.ZN(dbg_0_n_78_113), .A1(dbg_0_n_92), .A2(
      cpu_id[31]));
  NAND4_X1_LVT dbg_0_i_78_129 (.ZN(dbg_0_n_78_114), .A1(dbg_0_n_78_110), .A2(
      dbg_0_n_78_111), .A3(dbg_0_n_78_112), .A4(dbg_0_n_78_113));
  NAND2_X1_LVT dbg_0_i_49_7 (.ZN(dbg_0_n_49_7), .A1(dbg_0_n_49_2), .A2(
      dbg_0_n_49_6));
  NOR2_X1_LVT dbg_0_i_49_22 (.ZN(dbg_0_n_91), .A1(dbg_0_n_49_7), .A2(
      dbg_0_n_49_20));
  INV_X1_LVT dbg_0_i_49_18 (.ZN(dbg_0_n_49_18), .A(dbg_0_dbg_addr_in[5]));
  NAND2_X1_LVT dbg_0_i_49_17 (.ZN(dbg_0_n_49_17), .A1(dbg_0_dbg_addr_in[4]), .A2(
      dbg_0_n_49_18));
  INV_X1_LVT dbg_0_i_49_19 (.ZN(dbg_0_n_49_19), .A(dbg_0_n_49_17));
  NAND2_X1_LVT dbg_0_i_49_21 (.ZN(dbg_0_n_49_21), .A1(dbg_0_dbg_addr_in[3]), .A2(
      dbg_0_n_49_19));
  NOR2_X1_LVT dbg_0_i_49_30 (.ZN(dbg_0_n_99), .A1(dbg_0_n_49_7), .A2(
      dbg_0_n_49_21));
  AOI221_X1_LVT dbg_0_i_78_130 (.ZN(dbg_0_n_78_115), .A(dbg_0_n_78_114), .B1(
      dbg_0_n_91), .B2(cpu_id[15]), .C1(dbg_0_n_99), .C2(1'b0));
  INV_X1_LVT dbg_0_i_78_131 (.ZN(dbg_0_dbg_dout[15]), .A(dbg_0_n_78_115));
  NAND2_X1_LVT dbg_0_i_78_118 (.ZN(dbg_0_n_78_104), .A1(dbg_0_n_98), .A2(
      dbg_0_mem_cnt[14]));
  NAND2_X1_LVT dbg_0_i_78_119 (.ZN(dbg_0_n_78_105), .A1(dbg_0_n_96), .A2(
      dbg_mem_addr[14]));
  AND2_X1_LVT dbg_0_i_68_23 (.ZN(dbg_0_n_132), .A1(dbg_0_n_115), .A2(
      dbg_mem_din[14]));
  AOI222_X1_LVT dbg_0_i_71_28 (.ZN(dbg_0_n_71_14), .A1(dbg_0_mem_data_wr), .A2(
      dbg_0_dbg_din[14]), .B1(dbg_0_n_136), .B2(dbg_reg_din[14]), .C1(
      dbg_0_n_135), .C2(dbg_0_n_132));
  INV_X1_LVT dbg_0_i_71_29 (.ZN(dbg_0_n_151), .A(dbg_0_n_71_14));
  DFFR_X1_LVT \dbg_0_mem_data_reg[14] (.Q(dbg_0_mem_data[14]), .QN(), .CK(
      dbg_0_n_134), .D(dbg_0_n_151), .RN(dbg_0_n_104));
  NAND2_X1_LVT dbg_0_i_78_120 (.ZN(dbg_0_n_78_106), .A1(dbg_0_n_97), .A2(
      dbg_0_mem_data[14]));
  NAND2_X1_LVT dbg_0_i_78_121 (.ZN(dbg_0_n_78_107), .A1(dbg_0_n_92), .A2(
      cpu_id[30]));
  NAND4_X1_LVT dbg_0_i_78_122 (.ZN(dbg_0_n_78_108), .A1(dbg_0_n_78_104), .A2(
      dbg_0_n_78_105), .A3(dbg_0_n_78_106), .A4(dbg_0_n_78_107));
  AOI221_X1_LVT dbg_0_i_78_123 (.ZN(dbg_0_n_78_109), .A(dbg_0_n_78_108), .B1(
      dbg_0_n_91), .B2(cpu_id[14]), .C1(dbg_0_n_99), .C2(1'b0));
  INV_X1_LVT dbg_0_i_78_124 (.ZN(dbg_0_dbg_dout[14]), .A(dbg_0_n_78_109));
  NAND2_X1_LVT dbg_0_i_78_111 (.ZN(dbg_0_n_78_98), .A1(dbg_0_n_98), .A2(
      dbg_0_mem_cnt[13]));
  NAND2_X1_LVT dbg_0_i_78_112 (.ZN(dbg_0_n_78_99), .A1(dbg_0_n_96), .A2(
      dbg_mem_addr[13]));
  AND2_X1_LVT dbg_0_i_68_22 (.ZN(dbg_0_n_131), .A1(dbg_0_n_115), .A2(
      dbg_mem_din[13]));
  AOI222_X1_LVT dbg_0_i_71_26 (.ZN(dbg_0_n_71_13), .A1(dbg_0_mem_data_wr), .A2(
      dbg_0_dbg_din[13]), .B1(dbg_0_n_136), .B2(dbg_reg_din[13]), .C1(
      dbg_0_n_135), .C2(dbg_0_n_131));
  INV_X1_LVT dbg_0_i_71_27 (.ZN(dbg_0_n_150), .A(dbg_0_n_71_13));
  DFFR_X1_LVT \dbg_0_mem_data_reg[13] (.Q(dbg_0_mem_data[13]), .QN(), .CK(
      dbg_0_n_134), .D(dbg_0_n_150), .RN(dbg_0_n_104));
  NAND2_X1_LVT dbg_0_i_78_113 (.ZN(dbg_0_n_78_100), .A1(dbg_0_n_97), .A2(
      dbg_0_mem_data[13]));
  NAND2_X1_LVT dbg_0_i_78_114 (.ZN(dbg_0_n_78_101), .A1(dbg_0_n_92), .A2(
      cpu_id[29]));
  NAND4_X1_LVT dbg_0_i_78_115 (.ZN(dbg_0_n_78_102), .A1(dbg_0_n_78_98), .A2(
      dbg_0_n_78_99), .A3(dbg_0_n_78_100), .A4(dbg_0_n_78_101));
  AOI221_X1_LVT dbg_0_i_78_116 (.ZN(dbg_0_n_78_103), .A(dbg_0_n_78_102), .B1(
      dbg_0_n_91), .B2(cpu_id[13]), .C1(dbg_0_n_99), .C2(1'b0));
  INV_X1_LVT dbg_0_i_78_117 (.ZN(dbg_0_dbg_dout[13]), .A(dbg_0_n_78_103));
  NAND2_X1_LVT dbg_0_i_78_104 (.ZN(dbg_0_n_78_92), .A1(dbg_0_n_98), .A2(
      dbg_0_mem_cnt[12]));
  NAND2_X1_LVT dbg_0_i_78_105 (.ZN(dbg_0_n_78_93), .A1(dbg_0_n_96), .A2(
      dbg_mem_addr[12]));
  AND2_X1_LVT dbg_0_i_68_21 (.ZN(dbg_0_n_130), .A1(dbg_0_n_115), .A2(
      dbg_mem_din[12]));
  AOI222_X1_LVT dbg_0_i_71_24 (.ZN(dbg_0_n_71_12), .A1(dbg_0_mem_data_wr), .A2(
      dbg_0_dbg_din[12]), .B1(dbg_0_n_136), .B2(dbg_reg_din[12]), .C1(
      dbg_0_n_135), .C2(dbg_0_n_130));
  INV_X1_LVT dbg_0_i_71_25 (.ZN(dbg_0_n_149), .A(dbg_0_n_71_12));
  DFFR_X1_LVT \dbg_0_mem_data_reg[12] (.Q(dbg_0_mem_data[12]), .QN(), .CK(
      dbg_0_n_134), .D(dbg_0_n_149), .RN(dbg_0_n_104));
  NAND2_X1_LVT dbg_0_i_78_106 (.ZN(dbg_0_n_78_94), .A1(dbg_0_n_97), .A2(
      dbg_0_mem_data[12]));
  NAND2_X1_LVT dbg_0_i_78_107 (.ZN(dbg_0_n_78_95), .A1(dbg_0_n_92), .A2(
      cpu_id[28]));
  NAND4_X1_LVT dbg_0_i_78_108 (.ZN(dbg_0_n_78_96), .A1(dbg_0_n_78_92), .A2(
      dbg_0_n_78_93), .A3(dbg_0_n_78_94), .A4(dbg_0_n_78_95));
  AOI221_X1_LVT dbg_0_i_78_109 (.ZN(dbg_0_n_78_97), .A(dbg_0_n_78_96), .B1(
      dbg_0_n_91), .B2(cpu_id[12]), .C1(dbg_0_n_99), .C2(1'b0));
  INV_X1_LVT dbg_0_i_78_110 (.ZN(dbg_0_dbg_dout[12]), .A(dbg_0_n_78_97));
  NAND2_X1_LVT dbg_0_i_78_97 (.ZN(dbg_0_n_78_86), .A1(dbg_0_n_98), .A2(
      dbg_0_mem_cnt[11]));
  NAND2_X1_LVT dbg_0_i_78_98 (.ZN(dbg_0_n_78_87), .A1(dbg_0_n_96), .A2(
      dbg_mem_addr[11]));
  AND2_X1_LVT dbg_0_i_68_20 (.ZN(dbg_0_n_129), .A1(dbg_0_n_115), .A2(
      dbg_mem_din[11]));
  AOI222_X1_LVT dbg_0_i_71_22 (.ZN(dbg_0_n_71_11), .A1(dbg_0_mem_data_wr), .A2(
      dbg_0_dbg_din[11]), .B1(dbg_0_n_136), .B2(dbg_reg_din[11]), .C1(
      dbg_0_n_135), .C2(dbg_0_n_129));
  INV_X1_LVT dbg_0_i_71_23 (.ZN(dbg_0_n_148), .A(dbg_0_n_71_11));
  DFFR_X1_LVT \dbg_0_mem_data_reg[11] (.Q(dbg_0_mem_data[11]), .QN(), .CK(
      dbg_0_n_134), .D(dbg_0_n_148), .RN(dbg_0_n_104));
  NAND2_X1_LVT dbg_0_i_78_99 (.ZN(dbg_0_n_78_88), .A1(dbg_0_n_97), .A2(
      dbg_0_mem_data[11]));
  NAND2_X1_LVT dbg_0_i_78_100 (.ZN(dbg_0_n_78_89), .A1(dbg_0_n_92), .A2(
      cpu_id[27]));
  NAND4_X1_LVT dbg_0_i_78_101 (.ZN(dbg_0_n_78_90), .A1(dbg_0_n_78_86), .A2(
      dbg_0_n_78_87), .A3(dbg_0_n_78_88), .A4(dbg_0_n_78_89));
  AOI221_X1_LVT dbg_0_i_78_102 (.ZN(dbg_0_n_78_91), .A(dbg_0_n_78_90), .B1(
      dbg_0_n_91), .B2(cpu_id[11]), .C1(dbg_0_n_99), .C2(1'b0));
  INV_X1_LVT dbg_0_i_78_103 (.ZN(dbg_0_dbg_dout[11]), .A(dbg_0_n_78_91));
  NAND2_X1_LVT dbg_0_i_78_90 (.ZN(dbg_0_n_78_80), .A1(dbg_0_n_98), .A2(
      dbg_0_mem_cnt[10]));
  NAND2_X1_LVT dbg_0_i_78_91 (.ZN(dbg_0_n_78_81), .A1(dbg_0_n_96), .A2(
      dbg_mem_addr[10]));
  AND2_X1_LVT dbg_0_i_68_19 (.ZN(dbg_0_n_128), .A1(dbg_0_n_115), .A2(
      dbg_mem_din[10]));
  AOI222_X1_LVT dbg_0_i_71_20 (.ZN(dbg_0_n_71_10), .A1(dbg_0_mem_data_wr), .A2(
      dbg_0_dbg_din[10]), .B1(dbg_0_n_136), .B2(dbg_reg_din[10]), .C1(
      dbg_0_n_135), .C2(dbg_0_n_128));
  INV_X1_LVT dbg_0_i_71_21 (.ZN(dbg_0_n_147), .A(dbg_0_n_71_10));
  DFFR_X1_LVT \dbg_0_mem_data_reg[10] (.Q(dbg_0_mem_data[10]), .QN(), .CK(
      dbg_0_n_134), .D(dbg_0_n_147), .RN(dbg_0_n_104));
  NAND2_X1_LVT dbg_0_i_78_92 (.ZN(dbg_0_n_78_82), .A1(dbg_0_n_97), .A2(
      dbg_0_mem_data[10]));
  NAND2_X1_LVT dbg_0_i_78_93 (.ZN(dbg_0_n_78_83), .A1(dbg_0_n_92), .A2(
      cpu_id[26]));
  NAND4_X1_LVT dbg_0_i_78_94 (.ZN(dbg_0_n_78_84), .A1(dbg_0_n_78_80), .A2(
      dbg_0_n_78_81), .A3(dbg_0_n_78_82), .A4(dbg_0_n_78_83));
  AOI221_X1_LVT dbg_0_i_78_95 (.ZN(dbg_0_n_78_85), .A(dbg_0_n_78_84), .B1(
      dbg_0_n_91), .B2(cpu_id[10]), .C1(dbg_0_n_99), .C2(1'b0));
  INV_X1_LVT dbg_0_i_78_96 (.ZN(dbg_0_dbg_dout[10]), .A(dbg_0_n_78_85));
  NAND2_X1_LVT dbg_0_i_78_83 (.ZN(dbg_0_n_78_74), .A1(dbg_0_n_98), .A2(
      dbg_0_mem_cnt[9]));
  NAND2_X1_LVT dbg_0_i_78_84 (.ZN(dbg_0_n_78_75), .A1(dbg_0_n_96), .A2(
      dbg_mem_addr[9]));
  AND2_X1_LVT dbg_0_i_68_18 (.ZN(dbg_0_n_127), .A1(dbg_0_n_115), .A2(
      dbg_mem_din[9]));
  AOI222_X1_LVT dbg_0_i_71_18 (.ZN(dbg_0_n_71_9), .A1(dbg_0_mem_data_wr), .A2(
      dbg_0_dbg_din[9]), .B1(dbg_0_n_136), .B2(dbg_reg_din[9]), .C1(dbg_0_n_135), 
      .C2(dbg_0_n_127));
  INV_X1_LVT dbg_0_i_71_19 (.ZN(dbg_0_n_146), .A(dbg_0_n_71_9));
  DFFR_X1_LVT \dbg_0_mem_data_reg[9] (.Q(dbg_0_mem_data[9]), .QN(), .CK(
      dbg_0_n_134), .D(dbg_0_n_146), .RN(dbg_0_n_104));
  NAND2_X1_LVT dbg_0_i_78_85 (.ZN(dbg_0_n_78_76), .A1(dbg_0_n_97), .A2(
      dbg_0_mem_data[9]));
  NAND2_X1_LVT dbg_0_i_78_86 (.ZN(dbg_0_n_78_77), .A1(dbg_0_n_92), .A2(
      cpu_id[25]));
  NAND4_X1_LVT dbg_0_i_78_87 (.ZN(dbg_0_n_78_78), .A1(dbg_0_n_78_74), .A2(
      dbg_0_n_78_75), .A3(dbg_0_n_78_76), .A4(dbg_0_n_78_77));
  AOI221_X1_LVT dbg_0_i_78_88 (.ZN(dbg_0_n_78_79), .A(dbg_0_n_78_78), .B1(
      dbg_0_n_91), .B2(cpu_id[9]), .C1(dbg_0_n_99), .C2(1'b0));
  INV_X1_LVT dbg_0_i_78_89 (.ZN(dbg_0_dbg_dout[9]), .A(dbg_0_n_78_79));
  NAND2_X1_LVT dbg_0_i_78_76 (.ZN(dbg_0_n_78_68), .A1(dbg_0_n_98), .A2(
      dbg_0_mem_cnt[8]));
  NAND2_X1_LVT dbg_0_i_78_77 (.ZN(dbg_0_n_78_69), .A1(dbg_0_n_96), .A2(
      dbg_mem_addr[8]));
  AND2_X1_LVT dbg_0_i_68_17 (.ZN(dbg_0_n_126), .A1(dbg_mem_din[8]), .A2(
      dbg_0_n_115));
  AOI222_X1_LVT dbg_0_i_71_16 (.ZN(dbg_0_n_71_8), .A1(dbg_0_mem_data_wr), .A2(
      dbg_0_dbg_din[8]), .B1(dbg_0_n_136), .B2(dbg_reg_din[8]), .C1(dbg_0_n_135), 
      .C2(dbg_0_n_126));
  INV_X1_LVT dbg_0_i_71_17 (.ZN(dbg_0_n_145), .A(dbg_0_n_71_8));
  DFFR_X1_LVT \dbg_0_mem_data_reg[8] (.Q(dbg_0_mem_data[8]), .QN(), .CK(
      dbg_0_n_134), .D(dbg_0_n_145), .RN(dbg_0_n_104));
  NAND2_X1_LVT dbg_0_i_78_78 (.ZN(dbg_0_n_78_70), .A1(dbg_0_n_97), .A2(
      dbg_0_mem_data[8]));
  NAND2_X1_LVT dbg_0_i_78_79 (.ZN(dbg_0_n_78_71), .A1(dbg_0_n_92), .A2(
      cpu_id[24]));
  NAND4_X1_LVT dbg_0_i_78_80 (.ZN(dbg_0_n_78_72), .A1(dbg_0_n_78_68), .A2(
      dbg_0_n_78_69), .A3(dbg_0_n_78_70), .A4(dbg_0_n_78_71));
  AOI221_X1_LVT dbg_0_i_78_81 (.ZN(dbg_0_n_78_73), .A(dbg_0_n_78_72), .B1(
      dbg_0_n_91), .B2(cpu_id[8]), .C1(dbg_0_n_99), .C2(1'b0));
  INV_X1_LVT dbg_0_i_78_82 (.ZN(dbg_0_dbg_dout[8]), .A(dbg_0_n_78_73));
  NAND2_X1_LVT dbg_0_i_78_69 (.ZN(dbg_0_n_78_62), .A1(dbg_0_n_98), .A2(
      dbg_0_mem_cnt[7]));
  NAND2_X1_LVT dbg_0_i_78_70 (.ZN(dbg_0_n_78_63), .A1(dbg_0_n_96), .A2(
      dbg_mem_addr[7]));
  NOR2_X1_LVT dbg_0_i_67_1 (.ZN(dbg_0_n_116), .A1(dbg_0_n_115), .A2(
      dbg_mem_addr[0]));
  OR2_X1_LVT dbg_0_i_68_0 (.ZN(dbg_0_n_68_0), .A1(dbg_0_n_115), .A2(dbg_0_n_116));
  AND2_X1_LVT dbg_0_i_67_2 (.ZN(dbg_0_n_117), .A1(dbg_mem_addr[0]), .A2(
      dbg_0_mem_ctl[2]));
  AOI22_X1_LVT dbg_0_i_68_15 (.ZN(dbg_0_n_68_8), .A1(dbg_0_n_68_0), .A2(
      dbg_mem_din[7]), .B1(dbg_0_n_117), .B2(dbg_mem_din[15]));
  INV_X1_LVT dbg_0_i_68_16 (.ZN(dbg_0_n_125), .A(dbg_0_n_68_8));
  AOI222_X1_LVT dbg_0_i_71_14 (.ZN(dbg_0_n_71_7), .A1(dbg_0_mem_data_wr), .A2(
      dbg_0_dbg_din[7]), .B1(dbg_0_n_136), .B2(dbg_reg_din[7]), .C1(dbg_0_n_135), 
      .C2(dbg_0_n_125));
  INV_X1_LVT dbg_0_i_71_15 (.ZN(dbg_0_n_144), .A(dbg_0_n_71_7));
  DFFR_X1_LVT \dbg_0_mem_data_reg[7] (.Q(dbg_0_mem_data[7]), .QN(), .CK(
      dbg_0_n_134), .D(dbg_0_n_144), .RN(dbg_0_n_104));
  NAND2_X1_LVT dbg_0_i_78_71 (.ZN(dbg_0_n_78_64), .A1(dbg_0_n_97), .A2(
      dbg_0_mem_data[7]));
  NAND2_X1_LVT dbg_0_i_78_72 (.ZN(dbg_0_n_78_65), .A1(dbg_0_n_92), .A2(
      cpu_id[23]));
  NAND4_X1_LVT dbg_0_i_78_73 (.ZN(dbg_0_n_78_66), .A1(dbg_0_n_78_62), .A2(
      dbg_0_n_78_63), .A3(dbg_0_n_78_64), .A4(dbg_0_n_78_65));
  AOI221_X1_LVT dbg_0_i_78_74 (.ZN(dbg_0_n_78_67), .A(dbg_0_n_78_66), .B1(
      dbg_0_n_91), .B2(cpu_id[7]), .C1(dbg_0_n_99), .C2(1'b0));
  INV_X1_LVT dbg_0_i_78_75 (.ZN(dbg_0_dbg_dout[7]), .A(dbg_0_n_78_67));
  NAND2_X1_LVT dbg_0_i_78_60 (.ZN(dbg_0_n_78_54), .A1(dbg_0_n_96), .A2(
      dbg_mem_addr[6]));
  AOI22_X1_LVT dbg_0_i_68_13 (.ZN(dbg_0_n_68_7), .A1(dbg_0_n_68_0), .A2(
      dbg_mem_din[6]), .B1(dbg_0_n_117), .B2(dbg_mem_din[14]));
  INV_X1_LVT dbg_0_i_68_14 (.ZN(dbg_0_n_124), .A(dbg_0_n_68_7));
  AOI222_X1_LVT dbg_0_i_71_12 (.ZN(dbg_0_n_71_6), .A1(dbg_0_mem_data_wr), .A2(
      dbg_0_dbg_din[6]), .B1(dbg_0_n_136), .B2(dbg_reg_din[6]), .C1(dbg_0_n_135), 
      .C2(dbg_0_n_124));
  INV_X1_LVT dbg_0_i_71_13 (.ZN(dbg_0_n_143), .A(dbg_0_n_71_6));
  DFFR_X1_LVT \dbg_0_mem_data_reg[6] (.Q(dbg_0_mem_data[6]), .QN(), .CK(
      dbg_0_n_134), .D(dbg_0_n_143), .RN(dbg_0_n_104));
  NAND2_X1_LVT dbg_0_i_78_61 (.ZN(dbg_0_n_78_55), .A1(dbg_0_n_97), .A2(
      dbg_0_mem_data[6]));
  NAND2_X1_LVT dbg_0_i_49_9 (.ZN(dbg_0_n_49_9), .A1(dbg_0_n_49_4), .A2(
      dbg_0_n_49_6));
  NOR2_X1_LVT dbg_0_i_49_24 (.ZN(dbg_0_n_93), .A1(dbg_0_n_49_9), .A2(
      dbg_0_n_49_20));
  NAND2_X1_LVT dbg_0_i_78_62 (.ZN(dbg_0_n_78_56), .A1(dbg_0_n_93), .A2(
      dbg_cpu_reset));
  NAND2_X1_LVT dbg_0_i_78_63 (.ZN(dbg_0_n_78_57), .A1(dbg_0_n_92), .A2(
      cpu_id[22]));
  AND4_X1_LVT dbg_0_i_78_64 (.ZN(dbg_0_n_78_58), .A1(dbg_0_n_78_54), .A2(
      dbg_0_n_78_55), .A3(dbg_0_n_78_56), .A4(dbg_0_n_78_57));
  NAND2_X1_LVT dbg_0_i_78_65 (.ZN(dbg_0_n_78_59), .A1(dbg_0_n_91), .A2(cpu_id[6]));
  NAND2_X1_LVT dbg_0_i_78_66 (.ZN(dbg_0_n_78_60), .A1(dbg_0_n_99), .A2(1'b0));
  NAND2_X1_LVT dbg_0_i_78_67 (.ZN(dbg_0_n_78_61), .A1(dbg_0_n_98), .A2(
      dbg_0_mem_cnt[6]));
  NAND4_X1_LVT dbg_0_i_78_68 (.ZN(dbg_0_dbg_dout[6]), .A1(dbg_0_n_78_58), .A2(
      dbg_0_n_78_59), .A3(dbg_0_n_78_60), .A4(dbg_0_n_78_61));
  NAND2_X1_LVT dbg_0_i_78_51 (.ZN(dbg_0_n_78_46), .A1(dbg_0_n_96), .A2(
      dbg_mem_addr[5]));
  AOI22_X1_LVT dbg_0_i_68_11 (.ZN(dbg_0_n_68_6), .A1(dbg_0_n_68_0), .A2(
      dbg_mem_din[5]), .B1(dbg_0_n_117), .B2(dbg_mem_din[13]));
  INV_X1_LVT dbg_0_i_68_12 (.ZN(dbg_0_n_123), .A(dbg_0_n_68_6));
  AOI222_X1_LVT dbg_0_i_71_10 (.ZN(dbg_0_n_71_5), .A1(dbg_0_mem_data_wr), .A2(
      dbg_0_dbg_din[5]), .B1(dbg_0_n_136), .B2(dbg_reg_din[5]), .C1(dbg_0_n_135), 
      .C2(dbg_0_n_123));
  INV_X1_LVT dbg_0_i_71_11 (.ZN(dbg_0_n_142), .A(dbg_0_n_71_5));
  DFFR_X1_LVT \dbg_0_mem_data_reg[5] (.Q(dbg_0_mem_data[5]), .QN(), .CK(
      dbg_0_n_134), .D(dbg_0_n_142), .RN(dbg_0_n_104));
  NAND2_X1_LVT dbg_0_i_78_52 (.ZN(dbg_0_n_78_47), .A1(dbg_0_n_97), .A2(
      dbg_0_mem_data[5]));
  AND2_X1_LVT dbg_0_i_50_0 (.ZN(dbg_0_cpu_ctl_wr), .A1(dbg_0_dbg_wr), .A2(
      dbg_0_n_93));
  CLKGATETST_X1_LVT dbg_0_clk_gate_cpu_ctl_reg__0 (.GCK(dbg_0_n_105), .CK(
      dbg_clk), .E(dbg_0_cpu_ctl_wr), .SE(1'b0));
  DFFS_X1_LVT \dbg_0_cpu_ctl_reg[5] (.Q(dbg_0_cpu_ctl[2]), .QN(), .CK(
      dbg_0_n_105), .D(dbg_0_dbg_din[5]), .SN(dbg_0_n_104));
  NAND2_X1_LVT dbg_0_i_78_53 (.ZN(dbg_0_n_78_48), .A1(dbg_0_n_93), .A2(
      dbg_0_cpu_ctl[2]));
  NAND2_X1_LVT dbg_0_i_78_54 (.ZN(dbg_0_n_78_49), .A1(dbg_0_n_92), .A2(
      cpu_id[21]));
  AND4_X1_LVT dbg_0_i_78_55 (.ZN(dbg_0_n_78_50), .A1(dbg_0_n_78_46), .A2(
      dbg_0_n_78_47), .A3(dbg_0_n_78_48), .A4(dbg_0_n_78_49));
  NAND2_X1_LVT dbg_0_i_78_56 (.ZN(dbg_0_n_78_51), .A1(dbg_0_n_91), .A2(cpu_id[5]));
  NAND2_X1_LVT dbg_0_i_78_57 (.ZN(dbg_0_n_78_52), .A1(dbg_0_n_99), .A2(1'b0));
  NAND2_X1_LVT dbg_0_i_78_58 (.ZN(dbg_0_n_78_53), .A1(dbg_0_n_98), .A2(
      dbg_0_mem_cnt[5]));
  NAND4_X1_LVT dbg_0_i_78_59 (.ZN(dbg_0_dbg_dout[5]), .A1(dbg_0_n_78_50), .A2(
      dbg_0_n_78_51), .A3(dbg_0_n_78_52), .A4(dbg_0_n_78_53));
  NAND2_X1_LVT dbg_0_i_78_42 (.ZN(dbg_0_n_78_38), .A1(dbg_0_n_96), .A2(
      dbg_mem_addr[4]));
  AOI22_X1_LVT dbg_0_i_68_9 (.ZN(dbg_0_n_68_5), .A1(dbg_0_n_68_0), .A2(
      dbg_mem_din[4]), .B1(dbg_0_n_117), .B2(dbg_mem_din[12]));
  INV_X1_LVT dbg_0_i_68_10 (.ZN(dbg_0_n_122), .A(dbg_0_n_68_5));
  AOI222_X1_LVT dbg_0_i_71_8 (.ZN(dbg_0_n_71_4), .A1(dbg_0_mem_data_wr), .A2(
      dbg_0_dbg_din[4]), .B1(dbg_0_n_136), .B2(dbg_reg_din[4]), .C1(dbg_0_n_135), 
      .C2(dbg_0_n_122));
  INV_X1_LVT dbg_0_i_71_9 (.ZN(dbg_0_n_141), .A(dbg_0_n_71_4));
  DFFR_X1_LVT \dbg_0_mem_data_reg[4] (.Q(dbg_0_mem_data[4]), .QN(), .CK(
      dbg_0_n_134), .D(dbg_0_n_141), .RN(dbg_0_n_104));
  NAND2_X1_LVT dbg_0_i_78_43 (.ZN(dbg_0_n_78_39), .A1(dbg_0_n_97), .A2(
      dbg_0_mem_data[4]));
  CLKGATETST_X1_LVT dbg_0_clk_gate_cpu_ctl_reg__1 (.GCK(dbg_0_n_106), .CK(
      dbg_clk), .E(dbg_0_cpu_ctl_wr), .SE(1'b0));
  DFFS_X1_LVT \dbg_0_cpu_ctl_reg[4] (.Q(dbg_0_cpu_ctl[1]), .QN(), .CK(
      dbg_0_n_106), .D(dbg_0_dbg_din[4]), .SN(dbg_0_n_104));
  NAND2_X1_LVT dbg_0_i_78_44 (.ZN(dbg_0_n_78_40), .A1(dbg_0_n_93), .A2(
      dbg_0_cpu_ctl[1]));
  NAND2_X1_LVT dbg_0_i_78_45 (.ZN(dbg_0_n_78_41), .A1(dbg_0_n_92), .A2(
      cpu_id[20]));
  AND4_X1_LVT dbg_0_i_78_46 (.ZN(dbg_0_n_78_42), .A1(dbg_0_n_78_38), .A2(
      dbg_0_n_78_39), .A3(dbg_0_n_78_40), .A4(dbg_0_n_78_41));
  NAND2_X1_LVT dbg_0_i_78_47 (.ZN(dbg_0_n_78_43), .A1(dbg_0_n_91), .A2(cpu_id[4]));
  NAND2_X1_LVT dbg_0_i_78_48 (.ZN(dbg_0_n_78_44), .A1(dbg_0_n_99), .A2(1'b0));
  NAND2_X1_LVT dbg_0_i_78_49 (.ZN(dbg_0_n_78_45), .A1(dbg_0_n_98), .A2(
      dbg_0_mem_cnt[4]));
  NAND4_X1_LVT dbg_0_i_78_50 (.ZN(dbg_0_dbg_dout[4]), .A1(dbg_0_n_78_42), .A2(
      dbg_0_n_78_43), .A3(dbg_0_n_78_44), .A4(dbg_0_n_78_45));
  NAND2_X1_LVT dbg_0_i_78_29 (.ZN(dbg_0_n_78_26), .A1(dbg_0_n_99), .A2(1'b0));
  NAND2_X1_LVT dbg_0_i_78_30 (.ZN(dbg_0_n_78_27), .A1(dbg_0_n_98), .A2(
      dbg_0_mem_cnt[3]));
  NAND2_X1_LVT dbg_0_i_78_31 (.ZN(dbg_0_n_78_28), .A1(dbg_0_n_96), .A2(
      dbg_mem_addr[3]));
  AOI22_X1_LVT dbg_0_i_68_7 (.ZN(dbg_0_n_68_4), .A1(dbg_0_n_68_0), .A2(
      dbg_mem_din[3]), .B1(dbg_0_n_117), .B2(dbg_mem_din[11]));
  INV_X1_LVT dbg_0_i_68_8 (.ZN(dbg_0_n_121), .A(dbg_0_n_68_4));
  AOI222_X1_LVT dbg_0_i_71_6 (.ZN(dbg_0_n_71_3), .A1(dbg_0_mem_data_wr), .A2(
      dbg_0_dbg_din[3]), .B1(dbg_0_n_136), .B2(dbg_reg_din[3]), .C1(dbg_0_n_135), 
      .C2(dbg_0_n_121));
  INV_X1_LVT dbg_0_i_71_7 (.ZN(dbg_0_n_140), .A(dbg_0_n_71_3));
  DFFR_X1_LVT \dbg_0_mem_data_reg[3] (.Q(dbg_0_mem_data[3]), .QN(), .CK(
      dbg_0_n_134), .D(dbg_0_n_140), .RN(dbg_0_n_104));
  NAND2_X1_LVT dbg_0_i_78_32 (.ZN(dbg_0_n_78_29), .A1(dbg_0_n_97), .A2(
      dbg_0_mem_data[3]));
  NAND4_X1_LVT dbg_0_i_78_33 (.ZN(dbg_0_n_78_30), .A1(dbg_0_n_78_26), .A2(
      dbg_0_n_78_27), .A3(dbg_0_n_78_28), .A4(dbg_0_n_78_29));
  NAND2_X1_LVT dbg_0_i_78_34 (.ZN(dbg_0_n_78_31), .A1(dbg_0_n_95), .A2(
      dbg_0_mem_ctl[2]));
  NAND2_X1_LVT dbg_0_i_49_10 (.ZN(dbg_0_n_49_10), .A1(dbg_0_n_49_5), .A2(
      dbg_0_n_49_6));
  NOR2_X1_LVT dbg_0_i_49_25 (.ZN(dbg_0_n_94), .A1(dbg_0_n_49_10), .A2(
      dbg_0_n_49_20));
  NAND4_X1_LVT dbg_0_i_54_0 (.ZN(dbg_0_n_54_0), .A1(fe_mdb_in[0]), .A2(
      fe_mdb_in[1]), .A3(fe_mdb_in[6]), .A4(fe_mdb_in[8]));
  CLKGATETST_X1_LVT dbg_0_clk_gate_cpu_ctl_reg__2 (.GCK(dbg_0_n_107), .CK(
      dbg_clk), .E(dbg_0_cpu_ctl_wr), .SE(1'b0));
  DFFR_X1_LVT \dbg_0_cpu_ctl_reg[3] (.Q(dbg_0_cpu_ctl[0]), .QN(), .CK(dbg_0_n_107), 
      .D(dbg_0_dbg_din[3]), .RN(dbg_0_n_104));
  NAND4_X1_LVT dbg_0_i_54_1 (.ZN(dbg_0_n_54_1), .A1(fe_mdb_in[9]), .A2(
      fe_mdb_in[14]), .A3(dbg_0_cpu_ctl[0]), .A4(decode_noirq));
  NOR4_X1_LVT dbg_0_i_54_2 (.ZN(dbg_0_n_54_2), .A1(dbg_0_n_54_0), .A2(
      dbg_0_n_54_1), .A3(fe_mdb_in[13]), .A4(fe_mdb_in[15]));
  NOR4_X1_LVT dbg_0_i_54_3 (.ZN(dbg_0_n_54_3), .A1(fe_mdb_in[2]), .A2(
      fe_mdb_in[3]), .A3(fe_mdb_in[4]), .A4(fe_mdb_in[5]));
  NOR4_X1_LVT dbg_0_i_54_4 (.ZN(dbg_0_n_54_4), .A1(fe_mdb_in[7]), .A2(
      fe_mdb_in[10]), .A3(fe_mdb_in[11]), .A4(fe_mdb_in[12]));
  AND3_X1_LVT dbg_0_i_54_5 (.ZN(dbg_0_dbg_swbrk), .A1(dbg_0_n_54_2), .A2(
      dbg_0_n_54_3), .A3(dbg_0_n_54_4));
  INV_X1_LVT dbg_0_i_76_5 (.ZN(dbg_0_n_76_4), .A(dbg_0_dbg_din[3]));
  AOI21_X1_LVT dbg_0_i_76_6 (.ZN(dbg_0_n_76_5), .A(dbg_0_dbg_swbrk), .B1(
      dbg_0_n_76_4), .B2(dbg_0_cpu_stat[1]));
  AND2_X1_LVT dbg_0_i_50_1 (.ZN(dbg_0_n_100), .A1(dbg_0_dbg_wr), .A2(dbg_0_n_94));
  INV_X1_LVT dbg_0_i_76_2 (.ZN(dbg_0_n_76_2), .A(dbg_0_n_100));
  NOR2_X1_LVT dbg_0_i_76_7 (.ZN(dbg_0_n_76_6), .A1(dbg_0_cpu_stat[1]), .A2(
      dbg_0_dbg_swbrk));
  OAI22_X1_LVT dbg_0_i_76_8 (.ZN(dbg_0_n_155), .A1(dbg_0_n_76_5), .A2(
      dbg_0_n_76_2), .B1(dbg_0_n_76_6), .B2(dbg_0_n_100));
  DFFR_X1_LVT \dbg_0_cpu_stat_reg[3] (.Q(dbg_0_cpu_stat[1]), .QN(), .CK(dbg_clk), 
      .D(dbg_0_n_155), .RN(dbg_0_n_104));
  NAND2_X1_LVT dbg_0_i_78_35 (.ZN(dbg_0_n_78_32), .A1(dbg_0_n_94), .A2(
      dbg_0_cpu_stat[1]));
  NAND2_X1_LVT dbg_0_i_78_36 (.ZN(dbg_0_n_78_33), .A1(dbg_0_n_93), .A2(
      dbg_0_cpu_ctl[0]));
  NAND2_X1_LVT dbg_0_i_78_37 (.ZN(dbg_0_n_78_34), .A1(dbg_0_n_92), .A2(
      cpu_id[19]));
  NAND4_X1_LVT dbg_0_i_78_38 (.ZN(dbg_0_n_78_35), .A1(dbg_0_n_78_31), .A2(
      dbg_0_n_78_32), .A3(dbg_0_n_78_33), .A4(dbg_0_n_78_34));
  NOR2_X1_LVT dbg_0_i_78_39 (.ZN(dbg_0_n_78_36), .A1(dbg_0_n_78_30), .A2(
      dbg_0_n_78_35));
  NAND2_X1_LVT dbg_0_i_78_40 (.ZN(dbg_0_n_78_37), .A1(dbg_0_n_91), .A2(cpu_id[3]));
  NAND2_X1_LVT dbg_0_i_78_41 (.ZN(dbg_0_dbg_dout[3]), .A1(dbg_0_n_78_36), .A2(
      dbg_0_n_78_37));
  NAND2_X1_LVT dbg_0_i_78_18 (.ZN(dbg_0_n_78_16), .A1(dbg_0_n_91), .A2(cpu_id[2]));
  NAND2_X1_LVT dbg_0_i_78_19 (.ZN(dbg_0_n_78_17), .A1(dbg_0_n_99), .A2(1'b0));
  NAND2_X1_LVT dbg_0_i_78_20 (.ZN(dbg_0_n_78_18), .A1(dbg_0_n_98), .A2(
      dbg_0_mem_cnt[2]));
  NAND2_X1_LVT dbg_0_i_78_21 (.ZN(dbg_0_n_78_19), .A1(dbg_0_n_96), .A2(
      dbg_mem_addr[2]));
  NAND4_X1_LVT dbg_0_i_78_22 (.ZN(dbg_0_n_78_20), .A1(dbg_0_n_78_16), .A2(
      dbg_0_n_78_17), .A3(dbg_0_n_78_18), .A4(dbg_0_n_78_19));
  AOI22_X1_LVT dbg_0_i_68_5 (.ZN(dbg_0_n_68_3), .A1(dbg_0_n_68_0), .A2(
      dbg_mem_din[2]), .B1(dbg_0_n_117), .B2(dbg_mem_din[10]));
  INV_X1_LVT dbg_0_i_68_6 (.ZN(dbg_0_n_120), .A(dbg_0_n_68_3));
  AOI222_X1_LVT dbg_0_i_71_4 (.ZN(dbg_0_n_71_2), .A1(dbg_0_mem_data_wr), .A2(
      dbg_0_dbg_din[2]), .B1(dbg_0_n_136), .B2(dbg_reg_din[2]), .C1(dbg_0_n_135), 
      .C2(dbg_0_n_120));
  INV_X1_LVT dbg_0_i_71_5 (.ZN(dbg_0_n_139), .A(dbg_0_n_71_2));
  DFFR_X1_LVT \dbg_0_mem_data_reg[2] (.Q(dbg_0_mem_data[2]), .QN(), .CK(
      dbg_0_n_134), .D(dbg_0_n_139), .RN(dbg_0_n_104));
  NAND2_X1_LVT dbg_0_i_78_23 (.ZN(dbg_0_n_78_21), .A1(dbg_0_n_97), .A2(
      dbg_0_mem_data[2]));
  NAND2_X1_LVT dbg_0_i_78_24 (.ZN(dbg_0_n_78_22), .A1(dbg_0_n_95), .A2(
      dbg_0_mem_ctl[1]));
  INV_X1_LVT dbg_0_i_76_0 (.ZN(dbg_0_n_76_0), .A(dbg_0_dbg_din[2]));
  AOI21_X1_LVT dbg_0_i_76_1 (.ZN(dbg_0_n_76_1), .A(puc_pnd_set), .B1(
      dbg_0_n_76_0), .B2(dbg_0_cpu_stat[0]));
  NOR2_X1_LVT dbg_0_i_76_3 (.ZN(dbg_0_n_76_3), .A1(dbg_0_cpu_stat[0]), .A2(
      puc_pnd_set));
  OAI22_X1_LVT dbg_0_i_76_4 (.ZN(dbg_0_n_154), .A1(dbg_0_n_76_1), .A2(
      dbg_0_n_76_2), .B1(dbg_0_n_76_3), .B2(dbg_0_n_100));
  DFFR_X1_LVT \dbg_0_cpu_stat_reg[2] (.Q(dbg_0_cpu_stat[0]), .QN(), .CK(dbg_clk), 
      .D(dbg_0_n_154), .RN(dbg_0_n_104));
  NAND2_X1_LVT dbg_0_i_78_25 (.ZN(dbg_0_n_78_23), .A1(dbg_0_n_94), .A2(
      dbg_0_cpu_stat[0]));
  NAND2_X1_LVT dbg_0_i_78_26 (.ZN(dbg_0_n_78_24), .A1(dbg_0_n_92), .A2(
      cpu_id[18]));
  NAND4_X1_LVT dbg_0_i_78_27 (.ZN(dbg_0_n_78_25), .A1(dbg_0_n_78_21), .A2(
      dbg_0_n_78_22), .A3(dbg_0_n_78_23), .A4(dbg_0_n_78_24));
  OR2_X1_LVT dbg_0_i_78_28 (.ZN(dbg_0_dbg_dout[2]), .A1(dbg_0_n_78_20), .A2(
      dbg_0_n_78_25));
  NAND2_X1_LVT dbg_0_i_78_9 (.ZN(dbg_0_n_78_8), .A1(dbg_0_n_96), .A2(
      dbg_mem_addr[1]));
  AOI22_X1_LVT dbg_0_i_68_3 (.ZN(dbg_0_n_68_2), .A1(dbg_0_n_68_0), .A2(
      dbg_mem_din[1]), .B1(dbg_0_n_117), .B2(dbg_mem_din[9]));
  INV_X1_LVT dbg_0_i_68_4 (.ZN(dbg_0_n_119), .A(dbg_0_n_68_2));
  AOI222_X1_LVT dbg_0_i_71_2 (.ZN(dbg_0_n_71_1), .A1(dbg_0_mem_data_wr), .A2(
      dbg_0_dbg_din[1]), .B1(dbg_0_n_136), .B2(dbg_reg_din[1]), .C1(dbg_0_n_135), 
      .C2(dbg_0_n_119));
  INV_X1_LVT dbg_0_i_71_3 (.ZN(dbg_0_n_138), .A(dbg_0_n_71_1));
  DFFR_X1_LVT \dbg_0_mem_data_reg[1] (.Q(dbg_0_mem_data[1]), .QN(), .CK(
      dbg_0_n_134), .D(dbg_0_n_138), .RN(dbg_0_n_104));
  NAND2_X1_LVT dbg_0_i_78_10 (.ZN(dbg_0_n_78_9), .A1(dbg_0_n_97), .A2(
      dbg_0_mem_data[1]));
  NAND2_X1_LVT dbg_0_i_78_11 (.ZN(dbg_0_n_78_10), .A1(dbg_0_n_95), .A2(
      dbg_0_mem_ctl[0]));
  NAND2_X1_LVT dbg_0_i_78_12 (.ZN(dbg_0_n_78_11), .A1(dbg_0_n_92), .A2(
      cpu_id[17]));
  AND4_X1_LVT dbg_0_i_78_13 (.ZN(dbg_0_n_78_12), .A1(dbg_0_n_78_8), .A2(
      dbg_0_n_78_9), .A3(dbg_0_n_78_10), .A4(dbg_0_n_78_11));
  NAND2_X1_LVT dbg_0_i_78_14 (.ZN(dbg_0_n_78_13), .A1(dbg_0_n_91), .A2(cpu_id[1]));
  NAND2_X1_LVT dbg_0_i_78_15 (.ZN(dbg_0_n_78_14), .A1(dbg_0_n_99), .A2(1'b0));
  NAND2_X1_LVT dbg_0_i_78_16 (.ZN(dbg_0_n_78_15), .A1(dbg_0_n_98), .A2(
      dbg_0_mem_cnt[1]));
  NAND4_X1_LVT dbg_0_i_78_17 (.ZN(dbg_0_dbg_dout[1]), .A1(dbg_0_n_78_12), .A2(
      dbg_0_n_78_13), .A3(dbg_0_n_78_14), .A4(dbg_0_n_78_15));
  NAND2_X1_LVT dbg_0_i_78_0 (.ZN(dbg_0_n_78_0), .A1(dbg_mem_addr[0]), .A2(
      dbg_0_n_96));
  AOI22_X1_LVT dbg_0_i_68_1 (.ZN(dbg_0_n_68_1), .A1(dbg_0_n_68_0), .A2(
      dbg_mem_din[0]), .B1(dbg_mem_din[8]), .B2(dbg_0_n_117));
  INV_X1_LVT dbg_0_i_68_2 (.ZN(dbg_0_n_118), .A(dbg_0_n_68_1));
  AOI222_X1_LVT dbg_0_i_71_0 (.ZN(dbg_0_n_71_0), .A1(dbg_0_dbg_din[0]), .A2(
      dbg_0_mem_data_wr), .B1(dbg_reg_din[0]), .B2(dbg_0_n_136), .C1(dbg_0_n_118), 
      .C2(dbg_0_n_135));
  INV_X1_LVT dbg_0_i_71_1 (.ZN(dbg_0_n_137), .A(dbg_0_n_71_0));
  DFFR_X1_LVT \dbg_0_mem_data_reg[0] (.Q(dbg_0_mem_data[0]), .QN(), .CK(
      dbg_0_n_134), .D(dbg_0_n_137), .RN(dbg_0_n_104));
  NAND2_X1_LVT dbg_0_i_78_1 (.ZN(dbg_0_n_78_1), .A1(dbg_0_mem_data[0]), .A2(
      dbg_0_n_97));
  NAND2_X1_LVT dbg_0_i_78_2 (.ZN(dbg_0_n_78_2), .A1(cpu_halt_st), .A2(dbg_0_n_94));
  NAND2_X1_LVT dbg_0_i_78_3 (.ZN(dbg_0_n_78_3), .A1(cpu_id[16]), .A2(dbg_0_n_92));
  AND4_X1_LVT dbg_0_i_78_4 (.ZN(dbg_0_n_78_4), .A1(dbg_0_n_78_0), .A2(
      dbg_0_n_78_1), .A3(dbg_0_n_78_2), .A4(dbg_0_n_78_3));
  NAND2_X1_LVT dbg_0_i_78_5 (.ZN(dbg_0_n_78_5), .A1(cpu_id[0]), .A2(dbg_0_n_91));
  NAND2_X1_LVT dbg_0_i_78_6 (.ZN(dbg_0_n_78_6), .A1(1'b0), .A2(dbg_0_n_99));
  NAND2_X1_LVT dbg_0_i_78_7 (.ZN(dbg_0_n_78_7), .A1(dbg_0_mem_cnt[0]), .A2(
      dbg_0_n_98));
  NAND4_X1_LVT dbg_0_i_78_8 (.ZN(dbg_0_dbg_dout[0]), .A1(dbg_0_n_78_4), .A2(
      dbg_0_n_78_5), .A3(dbg_0_n_78_6), .A4(dbg_0_n_78_7));
  AND2_X1_LVT dbg_0_i_79_0 (.ZN(dbg_0_mem_burst_wr), .A1(dbg_0_mem_ctl[0]), .A2(
      dbg_0_mem_burst_start));
  INV_X1_LVT dbg_0_dbg_uart_0_i_4_0 (.ZN(dbg_0_dbg_uart_0_n_4_0), .A(
      dbg_0_dbg_rd_rdy));
  INV_X1_LVT dbg_0_dbg_uart_0_i_57_0 (.ZN(dbg_0_dbg_uart_0_n_136), .A(
      dbg_uart_rxd));
  INV_X1_LVT dbg_0_dbg_uart_0_sync_cell_uart_rxd_i_0_0 (.ZN(
      dbg_0_dbg_uart_0_sync_cell_uart_rxd_n_0), .A(dbg_rst));
  DFFR_X1_LVT \dbg_0_dbg_uart_0_sync_cell_uart_rxd_data_sync_reg[0] (.Q(
      dbg_0_dbg_uart_0_sync_cell_uart_rxd_n_1), .QN(), .CK(dbg_clk), .D(
      dbg_0_dbg_uart_0_n_136), .RN(dbg_0_dbg_uart_0_sync_cell_uart_rxd_n_0));
  DFFR_X1_LVT \dbg_0_dbg_uart_0_sync_cell_uart_rxd_data_sync_reg[1] (.Q(
      dbg_0_dbg_uart_0_uart_rxd_n), .QN(), .CK(dbg_clk), .D(
      dbg_0_dbg_uart_0_sync_cell_uart_rxd_n_1), .RN(
      dbg_0_dbg_uart_0_sync_cell_uart_rxd_n_0));
  INV_X1_LVT dbg_0_dbg_uart_0_i_0_0 (.ZN(dbg_0_dbg_uart_0_uart_rxd), .A(
      dbg_0_dbg_uart_0_uart_rxd_n));
  INV_X1_LVT dbg_0_dbg_uart_0_i_2_0 (.ZN(dbg_0_dbg_uart_0_n_2_0), .A(
      dbg_0_dbg_uart_0_uart_rxd));
  INV_X1_LVT dbg_0_dbg_uart_0_i_46_0 (.ZN(dbg_0_dbg_uart_0_n_130), .A(dbg_rst));
  DFFS_X1_LVT \dbg_0_dbg_uart_0_rxd_buf_reg[0] (.Q(dbg_0_dbg_uart_0_rxd_buf[0]), 
      .QN(), .CK(dbg_clk), .D(dbg_0_dbg_uart_0_uart_rxd), .SN(
      dbg_0_dbg_uart_0_n_130));
  INV_X1_LVT dbg_0_dbg_uart_0_i_2_1 (.ZN(dbg_0_dbg_uart_0_n_2_1), .A(
      dbg_0_dbg_uart_0_rxd_buf[0]));
  DFFS_X1_LVT \dbg_0_dbg_uart_0_rxd_buf_reg[1] (.Q(dbg_0_dbg_uart_0_rxd_buf[1]), 
      .QN(), .CK(dbg_clk), .D(dbg_0_dbg_uart_0_rxd_buf[0]), .SN(
      dbg_0_dbg_uart_0_n_130));
  INV_X1_LVT dbg_0_dbg_uart_0_i_2_2 (.ZN(dbg_0_dbg_uart_0_n_2_2), .A(
      dbg_0_dbg_uart_0_rxd_buf[1]));
  OAI222_X1_LVT dbg_0_dbg_uart_0_i_2_3 (.ZN(dbg_0_dbg_uart_0_rxd_maj_nxt), .A1(
      dbg_0_dbg_uart_0_n_2_0), .A2(dbg_0_dbg_uart_0_n_2_1), .B1(
      dbg_0_dbg_uart_0_n_2_1), .B2(dbg_0_dbg_uart_0_n_2_2), .C1(
      dbg_0_dbg_uart_0_n_2_0), .C2(dbg_0_dbg_uart_0_n_2_2));
  DFFS_X1_LVT dbg_0_dbg_uart_0_rxd_maj_reg (.Q(dbg_0_dbg_uart_0_rxd_maj), .QN(), 
      .CK(dbg_clk), .D(dbg_0_dbg_uart_0_rxd_maj_nxt), .SN(dbg_0_dbg_uart_0_n_130));
  INV_X1_LVT dbg_0_dbg_uart_0_i_4_36 (.ZN(dbg_0_dbg_uart_0_n_4_18), .A(
      dbg_0_dbg_uart_0_rxd_maj));
  NAND2_X1_LVT dbg_0_dbg_uart_0_i_4_37 (.ZN(dbg_0_dbg_uart_0_n_19), .A1(
      dbg_0_dbg_uart_0_n_4_18), .A2(dbg_0_dbg_uart_0_n_4_0));
  CLKGATETST_X1_LVT dbg_0_dbg_uart_0_clk_gate_sync_cnt_reg__16 (.GCK(
      dbg_0_dbg_uart_0_n_53), .CK(dbg_clk), .E(dbg_0_dbg_uart_0_n_76), .SE(1'b0));
  DFFR_X1_LVT \dbg_0_dbg_uart_0_sync_cnt_reg[1] (.Q(dbg_0_dbg_uart_0_n_54), .QN(), 
      .CK(dbg_0_dbg_uart_0_n_53), .D(dbg_0_dbg_uart_0_n_58), .RN(
      dbg_0_dbg_uart_0_n_130));
  INV_X1_LVT dbg_0_dbg_uart_0_i_21_0 (.ZN(dbg_0_dbg_uart_0_n_57), .A(
      dbg_0_dbg_uart_0_n_56));
  CLKGATETST_X1_LVT dbg_0_dbg_uart_0_clk_gate_sync_cnt_reg__17 (.GCK(
      dbg_0_dbg_uart_0_n_55), .CK(dbg_clk), .E(dbg_0_dbg_uart_0_n_76), .SE(1'b0));
  DFFR_X1_LVT \dbg_0_dbg_uart_0_sync_cnt_reg[0] (.Q(dbg_0_dbg_uart_0_n_56), .QN(), 
      .CK(dbg_0_dbg_uart_0_n_55), .D(dbg_0_dbg_uart_0_n_57), .RN(
      dbg_0_dbg_uart_0_n_130));
  HA_X1_LVT dbg_0_dbg_uart_0_i_21_1 (.CO(dbg_0_dbg_uart_0_n_21_0), .S(
      dbg_0_dbg_uart_0_n_58), .A(dbg_0_dbg_uart_0_n_54), .B(
      dbg_0_dbg_uart_0_n_56));
  HA_X1_LVT dbg_0_dbg_uart_0_i_21_2 (.CO(dbg_0_dbg_uart_0_n_21_1), .S(
      dbg_0_dbg_uart_0_n_59), .A(dbg_0_dbg_uart_0_n_52), .B(
      dbg_0_dbg_uart_0_n_21_0));
  CLKGATETST_X1_LVT dbg_0_dbg_uart_0_clk_gate_sync_cnt_reg__15 (.GCK(
      dbg_0_dbg_uart_0_n_51), .CK(dbg_clk), .E(dbg_0_dbg_uart_0_n_76), .SE(1'b0));
  DFFR_X1_LVT \dbg_0_dbg_uart_0_sync_cnt_reg[2] (.Q(dbg_0_dbg_uart_0_n_52), .QN(), 
      .CK(dbg_0_dbg_uart_0_n_51), .D(dbg_0_dbg_uart_0_n_59), .RN(
      dbg_0_dbg_uart_0_n_130));
  INV_X1_LVT dbg_0_dbg_uart_0_i_22_1 (.ZN(dbg_0_dbg_uart_0_n_22_1), .A(
      dbg_0_dbg_uart_0_n_52));
  NOR3_X1_LVT dbg_0_dbg_uart_0_i_8_4 (.ZN(dbg_0_dbg_uart_0_n_8_4), .A1(
      dbg_0_dbg_uart_0_n_8_3), .A2(dbg_0_dbg_uart_0_uart_state[0]), .A3(
      dbg_0_dbg_uart_0_uart_state[1]));
  INV_X1_LVT dbg_0_dbg_uart_0_i_8_5 (.ZN(dbg_0_dbg_uart_0_n_8_5), .A(
      dbg_0_dbg_uart_0_n_8_4));
  NAND3_X1_LVT dbg_0_dbg_uart_0_i_8_7 (.ZN(dbg_0_dbg_uart_0_n_8_7), .A1(
      dbg_0_dbg_uart_0_n_8_0), .A2(dbg_0_dbg_uart_0_uart_state[0]), .A3(
      dbg_0_dbg_uart_0_uart_state[2]));
  INV_X1_LVT dbg_0_dbg_uart_0_i_7_0 (.ZN(dbg_0_dbg_uart_0_n_7_0), .A(
      dbg_0_mem_burst));
  NOR2_X1_LVT dbg_0_dbg_uart_0_i_7_1 (.ZN(dbg_0_dbg_uart_0_n_22), .A1(
      dbg_0_dbg_uart_0_n_7_0), .A2(dbg_0_mem_burst_end));
  INV_X1_LVT dbg_0_dbg_uart_0_i_8_27 (.ZN(dbg_0_dbg_uart_0_n_8_26), .A(
      dbg_0_dbg_uart_0_n_22));
  INV_X1_LVT dbg_0_dbg_uart_0_i_8_20 (.ZN(dbg_0_dbg_uart_0_n_8_20), .A(
      dbg_0_mem_burst_wr));
  NAND2_X1_LVT dbg_0_dbg_uart_0_i_8_21 (.ZN(dbg_0_dbg_uart_0_n_8_21), .A1(
      dbg_0_dbg_uart_0_n_8_20), .A2(dbg_0_mem_burst_rd));
  INV_X1_LVT dbg_0_dbg_uart_0_i_8_29 (.ZN(dbg_0_dbg_uart_0_n_8_27), .A(
      dbg_0_dbg_uart_0_n_8_21));
  OR2_X1_LVT dbg_0_dbg_uart_0_i_8_15 (.ZN(dbg_0_dbg_uart_0_n_8_15), .A1(
      dbg_0_mem_burst_rd), .A2(dbg_0_mem_burst_wr));
  NOR2_X1_LVT dbg_0_dbg_uart_0_i_8_16 (.ZN(dbg_0_dbg_uart_0_n_8_16), .A1(
      dbg_0_dbg_uart_0_n_8_15), .A2(dbg_0_dbg_uart_0_xfer_buf[19]));
  AND2_X1_LVT dbg_0_dbg_uart_0_i_8_17 (.ZN(dbg_0_dbg_uart_0_n_8_17), .A1(
      dbg_0_dbg_uart_0_n_8_16), .A2(dbg_0_dbg_uart_0_xfer_buf[18]));
  INV_X1_LVT dbg_0_dbg_uart_0_i_8_30 (.ZN(dbg_0_dbg_uart_0_n_8_28), .A(
      dbg_0_dbg_uart_0_xfer_buf[18]));
  AOI211_X1_LVT dbg_0_dbg_uart_0_i_8_31 (.ZN(dbg_0_dbg_uart_0_n_8_29), .A(
      dbg_0_dbg_uart_0_n_8_27), .B(dbg_0_dbg_uart_0_n_8_17), .C1(
      dbg_0_dbg_uart_0_n_8_16), .C2(dbg_0_dbg_uart_0_n_8_28));
  INV_X1_LVT dbg_0_dbg_uart_0_i_8_24 (.ZN(dbg_0_dbg_uart_0_n_8_24), .A(
      dbg_0_dbg_uart_0_n_8_10));
  OAI221_X1_LVT dbg_0_dbg_uart_0_i_8_32 (.ZN(
      dbg_0_dbg_uart_0_uart_state_nxt_reg[2]), .A(dbg_0_dbg_uart_0_n_8_5), .B1(
      dbg_0_dbg_uart_0_n_8_7), .B2(dbg_0_dbg_uart_0_n_8_26), .C1(
      dbg_0_dbg_uart_0_n_8_29), .C2(dbg_0_dbg_uart_0_n_8_24));
  INV_X1_LVT dbg_0_dbg_uart_0_i_39_0 (.ZN(dbg_0_dbg_uart_0_n_119), .A(
      dbg_0_dbg_uart_0_xfer_bit[0]));
  AOI21_X1_LVT dbg_0_dbg_uart_0_i_41_1 (.ZN(dbg_0_dbg_uart_0_n_41_1), .A(
      dbg_0_dbg_uart_0_n_123), .B1(dbg_0_dbg_uart_0_n_41_0), .B2(
      dbg_0_dbg_uart_0_n_119));
  INV_X1_LVT dbg_0_dbg_uart_0_i_41_2 (.ZN(dbg_0_dbg_uart_0_n_124), .A(
      dbg_0_dbg_uart_0_n_41_1));
  INV_X1_LVT dbg_0_dbg_uart_0_i_42_0 (.ZN(dbg_0_dbg_uart_0_n_42_0), .A(
      dbg_0_dbg_uart_0_xfer_done));
  INV_X1_LVT dbg_0_dbg_uart_0_i_42_1 (.ZN(dbg_0_dbg_uart_0_n_42_1), .A(
      dbg_0_dbg_uart_0_n_123));
  NAND3_X1_LVT dbg_0_dbg_uart_0_i_42_2 (.ZN(dbg_0_dbg_uart_0_n_42_2), .A1(
      dbg_0_dbg_uart_0_n_42_0), .A2(dbg_0_dbg_uart_0_n_42_1), .A3(
      dbg_0_dbg_uart_0_xfer_bit_inc));
  NAND3_X1_LVT dbg_0_dbg_uart_0_i_42_3 (.ZN(dbg_0_dbg_uart_0_n_128), .A1(
      dbg_0_dbg_uart_0_n_42_2), .A2(dbg_0_dbg_uart_0_n_42_0), .A3(
      dbg_0_dbg_uart_0_n_42_1));
  CLKGATETST_X1_LVT dbg_0_dbg_uart_0_clk_gate_xfer_bit_reg (.GCK(
      dbg_0_dbg_uart_0_n_118), .CK(dbg_clk), .E(dbg_0_dbg_uart_0_n_128), .SE(
      1'b0));
  DFFR_X1_LVT \dbg_0_dbg_uart_0_xfer_bit_reg[0] (.Q(dbg_0_dbg_uart_0_xfer_bit[0]), 
      .QN(), .CK(dbg_0_dbg_uart_0_n_118), .D(dbg_0_dbg_uart_0_n_124), .RN(
      dbg_0_dbg_uart_0_n_130));
  HA_X1_LVT dbg_0_dbg_uart_0_i_39_1 (.CO(dbg_0_dbg_uart_0_n_39_0), .S(
      dbg_0_dbg_uart_0_n_120), .A(dbg_0_dbg_uart_0_xfer_bit[1]), .B(
      dbg_0_dbg_uart_0_xfer_bit[0]));
  AND2_X1_LVT dbg_0_dbg_uart_0_i_41_3 (.ZN(dbg_0_dbg_uart_0_n_125), .A1(
      dbg_0_dbg_uart_0_n_41_0), .A2(dbg_0_dbg_uart_0_n_120));
  DFFR_X1_LVT \dbg_0_dbg_uart_0_xfer_bit_reg[1] (.Q(dbg_0_dbg_uart_0_xfer_bit[1]), 
      .QN(), .CK(dbg_0_dbg_uart_0_n_118), .D(dbg_0_dbg_uart_0_n_125), .RN(
      dbg_0_dbg_uart_0_n_130));
  HA_X1_LVT dbg_0_dbg_uart_0_i_39_2 (.CO(dbg_0_dbg_uart_0_n_39_1), .S(
      dbg_0_dbg_uart_0_n_121), .A(dbg_0_dbg_uart_0_xfer_bit[2]), .B(
      dbg_0_dbg_uart_0_n_39_0));
  XNOR2_X1_LVT dbg_0_dbg_uart_0_i_39_3 (.ZN(dbg_0_dbg_uart_0_n_39_2), .A(
      dbg_0_dbg_uart_0_xfer_bit[3]), .B(dbg_0_dbg_uart_0_n_39_1));
  INV_X1_LVT dbg_0_dbg_uart_0_i_39_4 (.ZN(dbg_0_dbg_uart_0_n_122), .A(
      dbg_0_dbg_uart_0_n_39_2));
  AND2_X1_LVT dbg_0_dbg_uart_0_i_41_5 (.ZN(dbg_0_dbg_uart_0_n_127), .A1(
      dbg_0_dbg_uart_0_n_41_0), .A2(dbg_0_dbg_uart_0_n_122));
  DFFR_X1_LVT \dbg_0_dbg_uart_0_xfer_bit_reg[3] (.Q(dbg_0_dbg_uart_0_xfer_bit[3]), 
      .QN(), .CK(dbg_0_dbg_uart_0_n_118), .D(dbg_0_dbg_uart_0_n_127), .RN(
      dbg_0_dbg_uart_0_n_130));
  NOR4_X1_LVT dbg_0_dbg_uart_0_i_36_0 (.ZN(dbg_0_dbg_uart_0_n_116), .A1(
      dbg_0_dbg_uart_0_xfer_bit[0]), .A2(dbg_0_dbg_uart_0_xfer_bit[1]), .A3(
      dbg_0_dbg_uart_0_xfer_bit[2]), .A4(dbg_0_dbg_uart_0_xfer_bit[3]));
  OR3_X1_LVT dbg_0_dbg_uart_0_i_37_0 (.ZN(dbg_0_dbg_uart_0_n_117), .A1(
      dbg_0_dbg_uart_0_uart_state[0]), .A2(dbg_0_dbg_uart_0_uart_state[1]), .A3(
      dbg_0_dbg_uart_0_uart_state[2]));
  INV_X1_LVT dbg_0_dbg_uart_0_i_15_0 (.ZN(dbg_0_dbg_uart_0_n_15_0), .A(
      dbg_0_dbg_uart_0_rxd_maj));
  NOR2_X1_LVT dbg_0_dbg_uart_0_i_15_1 (.ZN(dbg_0_dbg_uart_0_rxd_fe), .A1(
      dbg_0_dbg_uart_0_n_15_0), .A2(dbg_0_dbg_uart_0_rxd_maj_nxt));
  AND3_X1_LVT dbg_0_dbg_uart_0_i_40_0 (.ZN(dbg_0_dbg_uart_0_n_40_0), .A1(
      dbg_0_dbg_uart_0_n_116), .A2(dbg_0_dbg_uart_0_n_117), .A3(
      dbg_0_dbg_uart_0_rxd_fe));
  INV_X1_LVT dbg_0_dbg_uart_0_i_13_5 (.ZN(dbg_0_dbg_uart_0_n_13_2), .A(
      dbg_0_dbg_uart_0_uart_state[2]));
  NOR3_X1_LVT dbg_0_dbg_uart_0_i_13_6 (.ZN(dbg_0_dbg_uart_0_n_28), .A1(
      dbg_0_dbg_uart_0_n_13_2), .A2(dbg_0_dbg_uart_0_uart_state[0]), .A3(
      dbg_0_dbg_uart_0_uart_state[1]));
  AOI21_X1_LVT dbg_0_dbg_uart_0_i_24_0 (.ZN(dbg_0_dbg_uart_0_n_24_0), .A(
      dbg_0_dbg_rd_rdy), .B1(dbg_0_dbg_uart_0_xfer_done), .B2(
      dbg_0_dbg_uart_0_n_28));
  INV_X1_LVT dbg_0_dbg_uart_0_i_24_1 (.ZN(dbg_0_dbg_uart_0_txd_start), .A(
      dbg_0_dbg_uart_0_n_24_0));
  OR2_X1_LVT dbg_0_dbg_uart_0_i_40_1 (.ZN(dbg_0_dbg_uart_0_n_123), .A1(
      dbg_0_dbg_uart_0_n_40_0), .A2(dbg_0_dbg_uart_0_txd_start));
  NOR2_X1_LVT dbg_0_dbg_uart_0_i_41_0 (.ZN(dbg_0_dbg_uart_0_n_41_0), .A1(
      dbg_0_dbg_uart_0_xfer_done), .A2(dbg_0_dbg_uart_0_n_123));
  AND2_X1_LVT dbg_0_dbg_uart_0_i_41_4 (.ZN(dbg_0_dbg_uart_0_n_126), .A1(
      dbg_0_dbg_uart_0_n_41_0), .A2(dbg_0_dbg_uart_0_n_121));
  DFFR_X1_LVT \dbg_0_dbg_uart_0_xfer_bit_reg[2] (.Q(dbg_0_dbg_uart_0_xfer_bit[2]), 
      .QN(), .CK(dbg_0_dbg_uart_0_n_118), .D(dbg_0_dbg_uart_0_n_126), .RN(
      dbg_0_dbg_uart_0_n_130));
  INV_X1_LVT dbg_0_dbg_uart_0_i_44_0 (.ZN(dbg_0_dbg_uart_0_n_44_0), .A(
      dbg_0_dbg_uart_0_xfer_bit[2]));
  INV_X1_LVT dbg_0_dbg_uart_0_i_13_0 (.ZN(dbg_0_dbg_uart_0_n_13_0), .A(
      dbg_0_dbg_uart_0_uart_state[1]));
  NOR3_X1_LVT dbg_0_dbg_uart_0_i_13_1 (.ZN(dbg_0_dbg_uart_0_n_25), .A1(
      dbg_0_dbg_uart_0_n_13_0), .A2(dbg_0_dbg_uart_0_uart_state[0]), .A3(
      dbg_0_dbg_uart_0_uart_state[2]));
  INV_X1_LVT dbg_0_dbg_uart_0_i_13_2 (.ZN(dbg_0_dbg_uart_0_n_13_1), .A(
      dbg_0_dbg_uart_0_uart_state[0]));
  NOR3_X1_LVT dbg_0_dbg_uart_0_i_13_4 (.ZN(dbg_0_dbg_uart_0_n_27), .A1(
      dbg_0_dbg_uart_0_n_13_1), .A2(dbg_0_dbg_uart_0_uart_state[1]), .A3(
      dbg_0_dbg_uart_0_uart_state[2]));
  NOR3_X1_LVT dbg_0_dbg_uart_0_i_13_3 (.ZN(dbg_0_dbg_uart_0_n_26), .A1(
      dbg_0_dbg_uart_0_n_13_0), .A2(dbg_0_dbg_uart_0_n_13_1), .A3(
      dbg_0_dbg_uart_0_uart_state[2]));
  OR3_X1_LVT dbg_0_dbg_uart_0_i_25_0 (.ZN(dbg_0_dbg_uart_0_rx_active), .A1(
      dbg_0_dbg_uart_0_n_25), .A2(dbg_0_dbg_uart_0_n_27), .A3(
      dbg_0_dbg_uart_0_n_26));
  NAND4_X1_LVT dbg_0_dbg_uart_0_i_44_1 (.ZN(dbg_0_dbg_uart_0_n_44_1), .A1(
      dbg_0_dbg_uart_0_n_44_0), .A2(dbg_0_dbg_uart_0_xfer_bit[1]), .A3(
      dbg_0_dbg_uart_0_xfer_bit[3]), .A4(dbg_0_dbg_uart_0_rx_active));
  INV_X1_LVT dbg_0_dbg_uart_0_i_44_2 (.ZN(dbg_0_dbg_uart_0_n_44_2), .A(
      dbg_0_dbg_uart_0_rx_active));
  NAND4_X1_LVT dbg_0_dbg_uart_0_i_44_3 (.ZN(dbg_0_dbg_uart_0_n_44_3), .A1(
      dbg_0_dbg_uart_0_n_44_2), .A2(dbg_0_dbg_uart_0_xfer_bit[0]), .A3(
      dbg_0_dbg_uart_0_xfer_bit[1]), .A4(dbg_0_dbg_uart_0_xfer_bit[3]));
  OAI22_X1_LVT dbg_0_dbg_uart_0_i_44_4 (.ZN(dbg_0_dbg_uart_0_xfer_done), .A1(
      dbg_0_dbg_uart_0_n_44_1), .A2(dbg_0_dbg_uart_0_xfer_bit[0]), .B1(
      dbg_0_dbg_uart_0_n_44_3), .B2(dbg_0_dbg_uart_0_xfer_bit[2]));
  NOR3_X1_LVT dbg_0_dbg_uart_0_i_11_0 (.ZN(dbg_0_dbg_uart_0_n_11_0), .A1(
      dbg_0_dbg_uart_0_xfer_done), .A2(dbg_0_mem_burst_rd), .A3(
      dbg_0_mem_burst_wr));
  NAND2_X1_LVT dbg_0_dbg_uart_0_i_14_0 (.ZN(dbg_0_dbg_uart_0_n_14_0), .A1(
      dbg_0_dbg_uart_0_n_29), .A2(dbg_0_dbg_uart_0_rxd_maj_nxt));
  NOR2_X1_LVT dbg_0_dbg_uart_0_i_14_1 (.ZN(dbg_0_dbg_uart_0_n_31), .A1(
      dbg_0_dbg_uart_0_n_14_0), .A2(dbg_0_dbg_uart_0_rxd_maj));
  NAND2_X1_LVT dbg_0_dbg_uart_0_i_11_1 (.ZN(dbg_0_dbg_uart_0_n_11_1), .A1(
      dbg_0_dbg_uart_0_n_31), .A2(dbg_0_dbg_uart_0_sync_busy));
  NAND2_X1_LVT dbg_0_dbg_uart_0_i_11_2 (.ZN(dbg_0_dbg_uart_0_n_24), .A1(
      dbg_0_dbg_uart_0_n_11_0), .A2(dbg_0_dbg_uart_0_n_11_1));
  CLKGATETST_X1_LVT dbg_0_dbg_uart_0_clk_gate_uart_state_reg (.GCK(
      dbg_0_dbg_uart_0_n_23), .CK(dbg_clk), .E(dbg_0_dbg_uart_0_n_24), .SE(1'b0));
  DFFR_X1_LVT \dbg_0_dbg_uart_0_uart_state_reg[2] (.Q(
      dbg_0_dbg_uart_0_uart_state[2]), .QN(), .CK(dbg_0_dbg_uart_0_n_23), .D(
      dbg_0_dbg_uart_0_uart_state_nxt_reg[2]), .RN(dbg_0_dbg_uart_0_n_130));
  INV_X1_LVT dbg_0_dbg_uart_0_i_8_3 (.ZN(dbg_0_dbg_uart_0_n_8_3), .A(
      dbg_0_dbg_uart_0_uart_state[2]));
  AND3_X1_LVT dbg_0_dbg_uart_0_i_8_10 (.ZN(dbg_0_dbg_uart_0_n_8_10), .A1(
      dbg_0_dbg_uart_0_n_8_0), .A2(dbg_0_dbg_uart_0_n_8_3), .A3(
      dbg_0_dbg_uart_0_uart_state[0]));
  INV_X1_LVT dbg_0_dbg_uart_0_i_8_18 (.ZN(dbg_0_dbg_uart_0_n_8_18), .A(
      dbg_0_dbg_uart_0_xfer_buf[19]));
  NOR2_X1_LVT dbg_0_dbg_uart_0_i_8_19 (.ZN(dbg_0_dbg_uart_0_n_8_19), .A1(
      dbg_0_dbg_uart_0_n_8_15), .A2(dbg_0_dbg_uart_0_n_8_18));
  OAI21_X1_LVT dbg_0_dbg_uart_0_i_8_26 (.ZN(dbg_0_dbg_uart_0_n_8_25), .A(
      dbg_0_dbg_uart_0_n_8_10), .B1(dbg_0_dbg_uart_0_n_8_19), .B2(
      dbg_0_mem_burst_wr));
  NAND3_X1_LVT dbg_0_dbg_uart_0_i_8_6 (.ZN(dbg_0_dbg_uart_0_n_8_6), .A1(
      dbg_0_dbg_uart_0_n_8_3), .A2(dbg_0_dbg_uart_0_uart_state[0]), .A3(
      dbg_0_dbg_uart_0_uart_state[1]));
  OAI211_X1_LVT dbg_0_dbg_uart_0_i_8_28 (.ZN(
      dbg_0_dbg_uart_0_uart_state_nxt_reg[1]), .A(dbg_0_dbg_uart_0_n_8_25), .B(
      dbg_0_dbg_uart_0_n_8_2), .C1(dbg_0_dbg_uart_0_n_8_6), .C2(
      dbg_0_dbg_uart_0_n_8_26));
  DFFR_X1_LVT \dbg_0_dbg_uart_0_uart_state_reg[1] (.Q(
      dbg_0_dbg_uart_0_uart_state[1]), .QN(), .CK(dbg_0_dbg_uart_0_n_23), .D(
      dbg_0_dbg_uart_0_uart_state_nxt_reg[1]), .RN(dbg_0_dbg_uart_0_n_130));
  INV_X1_LVT dbg_0_dbg_uart_0_i_8_0 (.ZN(dbg_0_dbg_uart_0_n_8_0), .A(
      dbg_0_dbg_uart_0_uart_state[1]));
  NOR3_X1_LVT dbg_0_dbg_uart_0_i_8_1 (.ZN(dbg_0_dbg_uart_0_n_8_1), .A1(
      dbg_0_dbg_uart_0_n_8_0), .A2(dbg_0_dbg_uart_0_uart_state[0]), .A3(
      dbg_0_dbg_uart_0_uart_state[2]));
  INV_X1_LVT dbg_0_dbg_uart_0_i_8_2 (.ZN(dbg_0_dbg_uart_0_n_8_2), .A(
      dbg_0_dbg_uart_0_n_8_1));
  NAND4_X1_LVT dbg_0_dbg_uart_0_i_8_8 (.ZN(dbg_0_dbg_uart_0_n_8_8), .A1(
      dbg_0_dbg_uart_0_n_8_2), .A2(dbg_0_dbg_uart_0_n_8_5), .A3(
      dbg_0_dbg_uart_0_n_8_6), .A4(dbg_0_dbg_uart_0_n_8_7));
  NOR3_X1_LVT dbg_0_dbg_uart_0_i_8_9 (.ZN(dbg_0_dbg_uart_0_n_8_9), .A1(
      dbg_0_dbg_uart_0_uart_state[0]), .A2(dbg_0_dbg_uart_0_uart_state[1]), .A3(
      dbg_0_dbg_uart_0_uart_state[2]));
  OR3_X1_LVT dbg_0_dbg_uart_0_i_8_11 (.ZN(dbg_0_dbg_uart_0_n_8_11), .A1(
      dbg_0_dbg_uart_0_n_8_8), .A2(dbg_0_dbg_uart_0_n_8_9), .A3(
      dbg_0_dbg_uart_0_n_8_10));
  NAND2_X1_LVT dbg_0_dbg_uart_0_i_8_12 (.ZN(dbg_0_dbg_uart_0_n_8_12), .A1(
      dbg_0_mem_ctl[2]), .A2(dbg_0_dbg_uart_0_n_22));
  AOI22_X1_LVT dbg_0_dbg_uart_0_i_8_13 (.ZN(dbg_0_dbg_uart_0_n_8_13), .A1(
      dbg_0_dbg_uart_0_n_8_6), .A2(dbg_0_dbg_uart_0_n_8_7), .B1(
      dbg_0_dbg_uart_0_n_8_12), .B2(dbg_0_dbg_uart_0_n_22));
  NOR4_X1_LVT dbg_0_dbg_uart_0_i_8_14 (.ZN(dbg_0_dbg_uart_0_n_8_14), .A1(
      dbg_0_dbg_uart_0_n_8_13), .A2(dbg_0_dbg_uart_0_n_8_4), .A3(
      dbg_0_dbg_uart_0_n_8_1), .A4(dbg_0_dbg_uart_0_n_8_9));
  NAND2_X1_LVT dbg_0_dbg_uart_0_i_8_22 (.ZN(dbg_0_dbg_uart_0_n_8_22), .A1(
      dbg_0_dbg_uart_0_n_8_21), .A2(dbg_0_dbg_uart_0_n_8_20));
  AOI221_X1_LVT dbg_0_dbg_uart_0_i_8_23 (.ZN(dbg_0_dbg_uart_0_n_8_23), .A(
      dbg_0_dbg_uart_0_n_8_17), .B1(dbg_0_dbg_uart_0_n_8_19), .B2(
      dbg_0_dbg_uart_0_xfer_buf[18]), .C1(dbg_0_dbg_uart_0_n_8_22), .C2(
      dbg_0_mem_ctl[2]));
  OAI211_X1_LVT dbg_0_dbg_uart_0_i_8_25 (.ZN(
      dbg_0_dbg_uart_0_uart_state_nxt_reg[0]), .A(dbg_0_dbg_uart_0_n_8_11), .B(
      dbg_0_dbg_uart_0_n_8_14), .C1(dbg_0_dbg_uart_0_n_8_23), .C2(
      dbg_0_dbg_uart_0_n_8_24));
  DFFR_X1_LVT \dbg_0_dbg_uart_0_uart_state_reg[0] (.Q(
      dbg_0_dbg_uart_0_uart_state[0]), .QN(), .CK(dbg_0_dbg_uart_0_n_23), .D(
      dbg_0_dbg_uart_0_uart_state_nxt_reg[0]), .RN(dbg_0_dbg_uart_0_n_130));
  NOR3_X1_LVT dbg_0_dbg_uart_0_i_13_7 (.ZN(dbg_0_dbg_uart_0_n_29), .A1(
      dbg_0_dbg_uart_0_uart_state[0]), .A2(dbg_0_dbg_uart_0_uart_state[1]), .A3(
      dbg_0_dbg_uart_0_uart_state[2]));
  AND2_X1_LVT dbg_0_dbg_uart_0_i_17_0 (.ZN(dbg_0_dbg_uart_0_n_33), .A1(
      dbg_0_dbg_uart_0_n_29), .A2(dbg_0_dbg_uart_0_rxd_fe));
  OR2_X1_LVT dbg_0_dbg_uart_0_i_18_0 (.ZN(dbg_0_dbg_uart_0_n_34), .A1(
      dbg_0_dbg_uart_0_n_31), .A2(dbg_0_dbg_uart_0_n_33));
  CLKGATETST_X1_LVT dbg_0_dbg_uart_0_clk_gate_sync_busy_reg (.GCK(
      dbg_0_dbg_uart_0_n_32), .CK(dbg_clk), .E(dbg_0_dbg_uart_0_n_34), .SE(1'b0));
  DFFR_X1_LVT dbg_0_dbg_uart_0_sync_busy_reg (.Q(dbg_0_dbg_uart_0_sync_busy), 
      .QN(), .CK(dbg_0_dbg_uart_0_n_32), .D(dbg_0_dbg_uart_0_n_33), .RN(
      dbg_0_dbg_uart_0_n_130));
  INV_X1_LVT dbg_0_dbg_uart_0_i_22_0 (.ZN(dbg_0_dbg_uart_0_n_22_0), .A(
      dbg_0_dbg_uart_0_sync_busy));
  NAND2_X1_LVT dbg_0_dbg_uart_0_i_22_2 (.ZN(dbg_0_dbg_uart_0_n_76), .A1(
      dbg_0_dbg_uart_0_n_22_1), .A2(dbg_0_dbg_uart_0_n_22_0));
  CLKGATETST_X1_LVT dbg_0_dbg_uart_0_clk_gate_sync_cnt_reg__14 (.GCK(
      dbg_0_dbg_uart_0_n_50), .CK(dbg_clk), .E(dbg_0_dbg_uart_0_n_76), .SE(1'b0));
  DFFS_X1_LVT \dbg_0_dbg_uart_0_sync_cnt_reg[3] (.Q(
      dbg_0_dbg_uart_0_bit_cnt_max[0]), .QN(), .CK(dbg_0_dbg_uart_0_n_50), .D(
      dbg_0_dbg_uart_0_n_60), .SN(dbg_0_dbg_uart_0_n_130));
  HA_X1_LVT dbg_0_dbg_uart_0_i_21_3 (.CO(dbg_0_dbg_uart_0_n_21_2), .S(
      dbg_0_dbg_uart_0_n_60), .A(dbg_0_dbg_uart_0_bit_cnt_max[0]), .B(
      dbg_0_dbg_uart_0_n_21_1));
  HA_X1_LVT dbg_0_dbg_uart_0_i_21_4 (.CO(dbg_0_dbg_uart_0_n_21_3), .S(
      dbg_0_dbg_uart_0_n_61), .A(dbg_0_dbg_uart_0_bit_cnt_max[1]), .B(
      dbg_0_dbg_uart_0_n_21_2));
  CLKGATETST_X1_LVT dbg_0_dbg_uart_0_clk_gate_sync_cnt_reg__13 (.GCK(
      dbg_0_dbg_uart_0_n_49), .CK(dbg_clk), .E(dbg_0_dbg_uart_0_n_76), .SE(1'b0));
  DFFS_X1_LVT \dbg_0_dbg_uart_0_sync_cnt_reg[4] (.Q(
      dbg_0_dbg_uart_0_bit_cnt_max[1]), .QN(), .CK(dbg_0_dbg_uart_0_n_49), .D(
      dbg_0_dbg_uart_0_n_61), .SN(dbg_0_dbg_uart_0_n_130));
  XOR2_X1_LVT dbg_0_dbg_uart_0_i_29_0 (.Z(dbg_0_dbg_uart_0_n_29_0), .A(
      dbg_0_dbg_uart_0_rxd_maj), .B(dbg_0_dbg_uart_0_rxd_maj_nxt));
  AND2_X1_LVT dbg_0_dbg_uart_0_i_29_1 (.ZN(dbg_0_dbg_uart_0_n_95), .A1(
      dbg_0_dbg_uart_0_n_29_0), .A2(dbg_0_dbg_uart_0_rx_active));
  OR2_X1_LVT dbg_0_dbg_uart_0_i_28_0 (.ZN(dbg_0_dbg_uart_0_n_94), .A1(
      dbg_0_dbg_uart_0_txd_start), .A2(dbg_0_dbg_uart_0_xfer_bit_inc));
  INV_X1_LVT dbg_0_dbg_uart_0_i_30_1 (.ZN(dbg_0_dbg_uart_0_n_30_0), .A(
      dbg_0_dbg_uart_0_n_94));
  NOR2_X1_LVT dbg_0_dbg_uart_0_i_30_2 (.ZN(dbg_0_dbg_uart_0_n_97), .A1(
      dbg_0_dbg_uart_0_n_30_0), .A2(dbg_0_dbg_uart_0_n_95));
  INV_X1_LVT dbg_0_dbg_uart_0_i_27_0 (.ZN(dbg_0_dbg_uart_0_n_78), .A(
      dbg_0_dbg_uart_0_xfer_cnt[0]));
  NOR2_X1_LVT dbg_0_dbg_uart_0_i_30_0 (.ZN(dbg_0_dbg_uart_0_n_96), .A1(
      dbg_0_dbg_uart_0_n_94), .A2(dbg_0_dbg_uart_0_n_95));
  AOI222_X1_LVT dbg_0_dbg_uart_0_i_31_0 (.ZN(dbg_0_dbg_uart_0_n_31_0), .A1(
      dbg_0_dbg_uart_0_bit_cnt_max[1]), .A2(dbg_0_dbg_uart_0_n_95), .B1(
      dbg_0_dbg_uart_0_bit_cnt_max[0]), .B2(dbg_0_dbg_uart_0_n_97), .C1(
      dbg_0_dbg_uart_0_n_78), .C2(dbg_0_dbg_uart_0_n_96));
  INV_X1_LVT dbg_0_dbg_uart_0_i_31_1 (.ZN(dbg_0_dbg_uart_0_n_98), .A(
      dbg_0_dbg_uart_0_n_31_0));
  INV_X1_LVT dbg_0_dbg_uart_0_i_33_0 (.ZN(dbg_0_dbg_uart_0_n_33_0), .A(
      dbg_0_dbg_uart_0_n_94));
  INV_X1_LVT dbg_0_dbg_uart_0_i_33_1 (.ZN(dbg_0_dbg_uart_0_n_33_1), .A(
      dbg_0_dbg_uart_0_n_95));
  XNOR2_X1_LVT dbg_0_dbg_uart_0_i_27_1 (.ZN(dbg_0_dbg_uart_0_n_79), .A(
      dbg_0_dbg_uart_0_xfer_cnt[1]), .B(dbg_0_dbg_uart_0_xfer_cnt[0]));
  NAND2_X1_LVT dbg_0_dbg_uart_0_i_31_2 (.ZN(dbg_0_dbg_uart_0_n_31_1), .A1(
      dbg_0_dbg_uart_0_n_96), .A2(dbg_0_dbg_uart_0_n_79));
  INV_X1_LVT dbg_0_dbg_uart_0_i_31_3 (.ZN(dbg_0_dbg_uart_0_n_31_2), .A(
      dbg_0_dbg_uart_0_n_95));
  HA_X1_LVT dbg_0_dbg_uart_0_i_21_5 (.CO(dbg_0_dbg_uart_0_n_21_4), .S(
      dbg_0_dbg_uart_0_n_62), .A(dbg_0_dbg_uart_0_bit_cnt_max[2]), .B(
      dbg_0_dbg_uart_0_n_21_3));
  CLKGATETST_X1_LVT dbg_0_dbg_uart_0_clk_gate_sync_cnt_reg__12 (.GCK(
      dbg_0_dbg_uart_0_n_48), .CK(dbg_clk), .E(dbg_0_dbg_uart_0_n_76), .SE(1'b0));
  DFFS_X1_LVT \dbg_0_dbg_uart_0_sync_cnt_reg[5] (.Q(
      dbg_0_dbg_uart_0_bit_cnt_max[2]), .QN(), .CK(dbg_0_dbg_uart_0_n_48), .D(
      dbg_0_dbg_uart_0_n_62), .SN(dbg_0_dbg_uart_0_n_130));
  INV_X1_LVT dbg_0_dbg_uart_0_i_31_4 (.ZN(dbg_0_dbg_uart_0_n_31_3), .A(
      dbg_0_dbg_uart_0_bit_cnt_max[2]));
  INV_X1_LVT dbg_0_dbg_uart_0_i_31_5 (.ZN(dbg_0_dbg_uart_0_n_31_4), .A(
      dbg_0_dbg_uart_0_bit_cnt_max[1]));
  INV_X1_LVT dbg_0_dbg_uart_0_i_31_6 (.ZN(dbg_0_dbg_uart_0_n_31_5), .A(
      dbg_0_dbg_uart_0_n_97));
  OAI221_X1_LVT dbg_0_dbg_uart_0_i_31_7 (.ZN(dbg_0_dbg_uart_0_n_99), .A(
      dbg_0_dbg_uart_0_n_31_1), .B1(dbg_0_dbg_uart_0_n_31_2), .B2(
      dbg_0_dbg_uart_0_n_31_3), .C1(dbg_0_dbg_uart_0_n_31_4), .C2(
      dbg_0_dbg_uart_0_n_31_5));
  DFFR_X1_LVT \dbg_0_dbg_uart_0_xfer_cnt_reg[1] (.Q(dbg_0_dbg_uart_0_xfer_cnt[1]), 
      .QN(), .CK(dbg_0_dbg_uart_0_n_77), .D(dbg_0_dbg_uart_0_n_99), .RN(
      dbg_0_dbg_uart_0_n_130));
  OR2_X1_LVT dbg_0_dbg_uart_0_i_27_2 (.ZN(dbg_0_dbg_uart_0_n_27_0), .A1(
      dbg_0_dbg_uart_0_xfer_cnt[1]), .A2(dbg_0_dbg_uart_0_xfer_cnt[0]));
  XNOR2_X1_LVT dbg_0_dbg_uart_0_i_27_3 (.ZN(dbg_0_dbg_uart_0_n_80), .A(
      dbg_0_dbg_uart_0_xfer_cnt[2]), .B(dbg_0_dbg_uart_0_n_27_0));
  NAND2_X1_LVT dbg_0_dbg_uart_0_i_31_8 (.ZN(dbg_0_dbg_uart_0_n_31_6), .A1(
      dbg_0_dbg_uart_0_n_96), .A2(dbg_0_dbg_uart_0_n_80));
  HA_X1_LVT dbg_0_dbg_uart_0_i_21_6 (.CO(dbg_0_dbg_uart_0_n_21_5), .S(
      dbg_0_dbg_uart_0_n_63), .A(dbg_0_dbg_uart_0_bit_cnt_max[3]), .B(
      dbg_0_dbg_uart_0_n_21_4));
  CLKGATETST_X1_LVT dbg_0_dbg_uart_0_clk_gate_sync_cnt_reg__11 (.GCK(
      dbg_0_dbg_uart_0_n_47), .CK(dbg_clk), .E(dbg_0_dbg_uart_0_n_76), .SE(1'b0));
  DFFS_X1_LVT \dbg_0_dbg_uart_0_sync_cnt_reg[6] (.Q(
      dbg_0_dbg_uart_0_bit_cnt_max[3]), .QN(), .CK(dbg_0_dbg_uart_0_n_47), .D(
      dbg_0_dbg_uart_0_n_63), .SN(dbg_0_dbg_uart_0_n_130));
  INV_X1_LVT dbg_0_dbg_uart_0_i_31_9 (.ZN(dbg_0_dbg_uart_0_n_31_7), .A(
      dbg_0_dbg_uart_0_bit_cnt_max[3]));
  OAI221_X1_LVT dbg_0_dbg_uart_0_i_31_10 (.ZN(dbg_0_dbg_uart_0_n_100), .A(
      dbg_0_dbg_uart_0_n_31_6), .B1(dbg_0_dbg_uart_0_n_31_2), .B2(
      dbg_0_dbg_uart_0_n_31_7), .C1(dbg_0_dbg_uart_0_n_31_5), .C2(
      dbg_0_dbg_uart_0_n_31_3));
  DFFR_X1_LVT \dbg_0_dbg_uart_0_xfer_cnt_reg[2] (.Q(dbg_0_dbg_uart_0_xfer_cnt[2]), 
      .QN(), .CK(dbg_0_dbg_uart_0_n_77), .D(dbg_0_dbg_uart_0_n_100), .RN(
      dbg_0_dbg_uart_0_n_130));
  OR2_X1_LVT dbg_0_dbg_uart_0_i_27_4 (.ZN(dbg_0_dbg_uart_0_n_27_1), .A1(
      dbg_0_dbg_uart_0_xfer_cnt[2]), .A2(dbg_0_dbg_uart_0_n_27_0));
  XNOR2_X1_LVT dbg_0_dbg_uart_0_i_27_5 (.ZN(dbg_0_dbg_uart_0_n_81), .A(
      dbg_0_dbg_uart_0_xfer_cnt[3]), .B(dbg_0_dbg_uart_0_n_27_1));
  NAND2_X1_LVT dbg_0_dbg_uart_0_i_31_11 (.ZN(dbg_0_dbg_uart_0_n_31_8), .A1(
      dbg_0_dbg_uart_0_n_96), .A2(dbg_0_dbg_uart_0_n_81));
  HA_X1_LVT dbg_0_dbg_uart_0_i_21_7 (.CO(dbg_0_dbg_uart_0_n_21_6), .S(
      dbg_0_dbg_uart_0_n_64), .A(dbg_0_dbg_uart_0_bit_cnt_max[4]), .B(
      dbg_0_dbg_uart_0_n_21_5));
  CLKGATETST_X1_LVT dbg_0_dbg_uart_0_clk_gate_sync_cnt_reg__10 (.GCK(
      dbg_0_dbg_uart_0_n_46), .CK(dbg_clk), .E(dbg_0_dbg_uart_0_n_76), .SE(1'b0));
  DFFS_X1_LVT \dbg_0_dbg_uart_0_sync_cnt_reg[7] (.Q(
      dbg_0_dbg_uart_0_bit_cnt_max[4]), .QN(), .CK(dbg_0_dbg_uart_0_n_46), .D(
      dbg_0_dbg_uart_0_n_64), .SN(dbg_0_dbg_uart_0_n_130));
  INV_X1_LVT dbg_0_dbg_uart_0_i_31_12 (.ZN(dbg_0_dbg_uart_0_n_31_9), .A(
      dbg_0_dbg_uart_0_bit_cnt_max[4]));
  OAI221_X1_LVT dbg_0_dbg_uart_0_i_31_13 (.ZN(dbg_0_dbg_uart_0_n_101), .A(
      dbg_0_dbg_uart_0_n_31_8), .B1(dbg_0_dbg_uart_0_n_31_2), .B2(
      dbg_0_dbg_uart_0_n_31_9), .C1(dbg_0_dbg_uart_0_n_31_5), .C2(
      dbg_0_dbg_uart_0_n_31_7));
  DFFR_X1_LVT \dbg_0_dbg_uart_0_xfer_cnt_reg[3] (.Q(dbg_0_dbg_uart_0_xfer_cnt[3]), 
      .QN(), .CK(dbg_0_dbg_uart_0_n_77), .D(dbg_0_dbg_uart_0_n_101), .RN(
      dbg_0_dbg_uart_0_n_130));
  NOR4_X1_LVT dbg_0_dbg_uart_0_i_32_0 (.ZN(dbg_0_dbg_uart_0_n_32_0), .A1(
      dbg_0_dbg_uart_0_xfer_cnt[0]), .A2(dbg_0_dbg_uart_0_xfer_cnt[1]), .A3(
      dbg_0_dbg_uart_0_xfer_cnt[2]), .A4(dbg_0_dbg_uart_0_xfer_cnt[3]));
  OR2_X1_LVT dbg_0_dbg_uart_0_i_27_6 (.ZN(dbg_0_dbg_uart_0_n_27_2), .A1(
      dbg_0_dbg_uart_0_xfer_cnt[3]), .A2(dbg_0_dbg_uart_0_n_27_1));
  XNOR2_X1_LVT dbg_0_dbg_uart_0_i_27_7 (.ZN(dbg_0_dbg_uart_0_n_82), .A(
      dbg_0_dbg_uart_0_xfer_cnt[4]), .B(dbg_0_dbg_uart_0_n_27_2));
  NAND2_X1_LVT dbg_0_dbg_uart_0_i_31_14 (.ZN(dbg_0_dbg_uart_0_n_31_10), .A1(
      dbg_0_dbg_uart_0_n_96), .A2(dbg_0_dbg_uart_0_n_82));
  HA_X1_LVT dbg_0_dbg_uart_0_i_21_8 (.CO(dbg_0_dbg_uart_0_n_21_7), .S(
      dbg_0_dbg_uart_0_n_65), .A(dbg_0_dbg_uart_0_bit_cnt_max[5]), .B(
      dbg_0_dbg_uart_0_n_21_6));
  CLKGATETST_X1_LVT dbg_0_dbg_uart_0_clk_gate_sync_cnt_reg__9 (.GCK(
      dbg_0_dbg_uart_0_n_45), .CK(dbg_clk), .E(dbg_0_dbg_uart_0_n_76), .SE(1'b0));
  DFFS_X1_LVT \dbg_0_dbg_uart_0_sync_cnt_reg[8] (.Q(
      dbg_0_dbg_uart_0_bit_cnt_max[5]), .QN(), .CK(dbg_0_dbg_uart_0_n_45), .D(
      dbg_0_dbg_uart_0_n_65), .SN(dbg_0_dbg_uart_0_n_130));
  INV_X1_LVT dbg_0_dbg_uart_0_i_31_15 (.ZN(dbg_0_dbg_uart_0_n_31_11), .A(
      dbg_0_dbg_uart_0_bit_cnt_max[5]));
  OAI221_X1_LVT dbg_0_dbg_uart_0_i_31_16 (.ZN(dbg_0_dbg_uart_0_n_102), .A(
      dbg_0_dbg_uart_0_n_31_10), .B1(dbg_0_dbg_uart_0_n_31_2), .B2(
      dbg_0_dbg_uart_0_n_31_11), .C1(dbg_0_dbg_uart_0_n_31_5), .C2(
      dbg_0_dbg_uart_0_n_31_9));
  DFFR_X1_LVT \dbg_0_dbg_uart_0_xfer_cnt_reg[4] (.Q(dbg_0_dbg_uart_0_xfer_cnt[4]), 
      .QN(), .CK(dbg_0_dbg_uart_0_n_77), .D(dbg_0_dbg_uart_0_n_102), .RN(
      dbg_0_dbg_uart_0_n_130));
  OR2_X1_LVT dbg_0_dbg_uart_0_i_27_8 (.ZN(dbg_0_dbg_uart_0_n_27_3), .A1(
      dbg_0_dbg_uart_0_xfer_cnt[4]), .A2(dbg_0_dbg_uart_0_n_27_2));
  XNOR2_X1_LVT dbg_0_dbg_uart_0_i_27_9 (.ZN(dbg_0_dbg_uart_0_n_83), .A(
      dbg_0_dbg_uart_0_xfer_cnt[5]), .B(dbg_0_dbg_uart_0_n_27_3));
  NAND2_X1_LVT dbg_0_dbg_uart_0_i_31_17 (.ZN(dbg_0_dbg_uart_0_n_31_12), .A1(
      dbg_0_dbg_uart_0_n_96), .A2(dbg_0_dbg_uart_0_n_83));
  HA_X1_LVT dbg_0_dbg_uart_0_i_21_9 (.CO(dbg_0_dbg_uart_0_n_21_8), .S(
      dbg_0_dbg_uart_0_n_66), .A(dbg_0_dbg_uart_0_bit_cnt_max[6]), .B(
      dbg_0_dbg_uart_0_n_21_7));
  CLKGATETST_X1_LVT dbg_0_dbg_uart_0_clk_gate_sync_cnt_reg__8 (.GCK(
      dbg_0_dbg_uart_0_n_44), .CK(dbg_clk), .E(dbg_0_dbg_uart_0_n_76), .SE(1'b0));
  DFFS_X1_LVT \dbg_0_dbg_uart_0_sync_cnt_reg[9] (.Q(
      dbg_0_dbg_uart_0_bit_cnt_max[6]), .QN(), .CK(dbg_0_dbg_uart_0_n_44), .D(
      dbg_0_dbg_uart_0_n_66), .SN(dbg_0_dbg_uart_0_n_130));
  INV_X1_LVT dbg_0_dbg_uart_0_i_31_18 (.ZN(dbg_0_dbg_uart_0_n_31_13), .A(
      dbg_0_dbg_uart_0_bit_cnt_max[6]));
  OAI221_X1_LVT dbg_0_dbg_uart_0_i_31_19 (.ZN(dbg_0_dbg_uart_0_n_103), .A(
      dbg_0_dbg_uart_0_n_31_12), .B1(dbg_0_dbg_uart_0_n_31_2), .B2(
      dbg_0_dbg_uart_0_n_31_13), .C1(dbg_0_dbg_uart_0_n_31_5), .C2(
      dbg_0_dbg_uart_0_n_31_11));
  DFFR_X1_LVT \dbg_0_dbg_uart_0_xfer_cnt_reg[5] (.Q(dbg_0_dbg_uart_0_xfer_cnt[5]), 
      .QN(), .CK(dbg_0_dbg_uart_0_n_77), .D(dbg_0_dbg_uart_0_n_103), .RN(
      dbg_0_dbg_uart_0_n_130));
  OR2_X1_LVT dbg_0_dbg_uart_0_i_27_10 (.ZN(dbg_0_dbg_uart_0_n_27_4), .A1(
      dbg_0_dbg_uart_0_xfer_cnt[5]), .A2(dbg_0_dbg_uart_0_n_27_3));
  XNOR2_X1_LVT dbg_0_dbg_uart_0_i_27_11 (.ZN(dbg_0_dbg_uart_0_n_84), .A(
      dbg_0_dbg_uart_0_xfer_cnt[6]), .B(dbg_0_dbg_uart_0_n_27_4));
  NAND2_X1_LVT dbg_0_dbg_uart_0_i_31_20 (.ZN(dbg_0_dbg_uart_0_n_31_14), .A1(
      dbg_0_dbg_uart_0_n_96), .A2(dbg_0_dbg_uart_0_n_84));
  HA_X1_LVT dbg_0_dbg_uart_0_i_21_10 (.CO(dbg_0_dbg_uart_0_n_21_9), .S(
      dbg_0_dbg_uart_0_n_67), .A(dbg_0_dbg_uart_0_bit_cnt_max[7]), .B(
      dbg_0_dbg_uart_0_n_21_8));
  CLKGATETST_X1_LVT dbg_0_dbg_uart_0_clk_gate_sync_cnt_reg__7 (.GCK(
      dbg_0_dbg_uart_0_n_43), .CK(dbg_clk), .E(dbg_0_dbg_uart_0_n_76), .SE(1'b0));
  DFFS_X1_LVT \dbg_0_dbg_uart_0_sync_cnt_reg[10] (.Q(
      dbg_0_dbg_uart_0_bit_cnt_max[7]), .QN(), .CK(dbg_0_dbg_uart_0_n_43), .D(
      dbg_0_dbg_uart_0_n_67), .SN(dbg_0_dbg_uart_0_n_130));
  INV_X1_LVT dbg_0_dbg_uart_0_i_31_21 (.ZN(dbg_0_dbg_uart_0_n_31_15), .A(
      dbg_0_dbg_uart_0_bit_cnt_max[7]));
  OAI221_X1_LVT dbg_0_dbg_uart_0_i_31_22 (.ZN(dbg_0_dbg_uart_0_n_104), .A(
      dbg_0_dbg_uart_0_n_31_14), .B1(dbg_0_dbg_uart_0_n_31_2), .B2(
      dbg_0_dbg_uart_0_n_31_15), .C1(dbg_0_dbg_uart_0_n_31_5), .C2(
      dbg_0_dbg_uart_0_n_31_13));
  DFFR_X1_LVT \dbg_0_dbg_uart_0_xfer_cnt_reg[6] (.Q(dbg_0_dbg_uart_0_xfer_cnt[6]), 
      .QN(), .CK(dbg_0_dbg_uart_0_n_77), .D(dbg_0_dbg_uart_0_n_104), .RN(
      dbg_0_dbg_uart_0_n_130));
  OR2_X1_LVT dbg_0_dbg_uart_0_i_27_12 (.ZN(dbg_0_dbg_uart_0_n_27_5), .A1(
      dbg_0_dbg_uart_0_xfer_cnt[6]), .A2(dbg_0_dbg_uart_0_n_27_4));
  XNOR2_X1_LVT dbg_0_dbg_uart_0_i_27_13 (.ZN(dbg_0_dbg_uart_0_n_85), .A(
      dbg_0_dbg_uart_0_xfer_cnt[7]), .B(dbg_0_dbg_uart_0_n_27_5));
  NAND2_X1_LVT dbg_0_dbg_uart_0_i_31_23 (.ZN(dbg_0_dbg_uart_0_n_31_16), .A1(
      dbg_0_dbg_uart_0_n_96), .A2(dbg_0_dbg_uart_0_n_85));
  HA_X1_LVT dbg_0_dbg_uart_0_i_21_11 (.CO(dbg_0_dbg_uart_0_n_21_10), .S(
      dbg_0_dbg_uart_0_n_68), .A(dbg_0_dbg_uart_0_bit_cnt_max[8]), .B(
      dbg_0_dbg_uart_0_n_21_9));
  CLKGATETST_X1_LVT dbg_0_dbg_uart_0_clk_gate_sync_cnt_reg__6 (.GCK(
      dbg_0_dbg_uart_0_n_42), .CK(dbg_clk), .E(dbg_0_dbg_uart_0_n_76), .SE(1'b0));
  DFFS_X1_LVT \dbg_0_dbg_uart_0_sync_cnt_reg[11] (.Q(
      dbg_0_dbg_uart_0_bit_cnt_max[8]), .QN(), .CK(dbg_0_dbg_uart_0_n_42), .D(
      dbg_0_dbg_uart_0_n_68), .SN(dbg_0_dbg_uart_0_n_130));
  INV_X1_LVT dbg_0_dbg_uart_0_i_31_24 (.ZN(dbg_0_dbg_uart_0_n_31_17), .A(
      dbg_0_dbg_uart_0_bit_cnt_max[8]));
  OAI221_X1_LVT dbg_0_dbg_uart_0_i_31_25 (.ZN(dbg_0_dbg_uart_0_n_105), .A(
      dbg_0_dbg_uart_0_n_31_16), .B1(dbg_0_dbg_uart_0_n_31_2), .B2(
      dbg_0_dbg_uart_0_n_31_17), .C1(dbg_0_dbg_uart_0_n_31_5), .C2(
      dbg_0_dbg_uart_0_n_31_15));
  DFFR_X1_LVT \dbg_0_dbg_uart_0_xfer_cnt_reg[7] (.Q(dbg_0_dbg_uart_0_xfer_cnt[7]), 
      .QN(), .CK(dbg_0_dbg_uart_0_n_77), .D(dbg_0_dbg_uart_0_n_105), .RN(
      dbg_0_dbg_uart_0_n_130));
  NOR4_X1_LVT dbg_0_dbg_uart_0_i_32_1 (.ZN(dbg_0_dbg_uart_0_n_32_1), .A1(
      dbg_0_dbg_uart_0_xfer_cnt[4]), .A2(dbg_0_dbg_uart_0_xfer_cnt[5]), .A3(
      dbg_0_dbg_uart_0_xfer_cnt[6]), .A4(dbg_0_dbg_uart_0_xfer_cnt[7]));
  OR2_X1_LVT dbg_0_dbg_uart_0_i_27_14 (.ZN(dbg_0_dbg_uart_0_n_27_6), .A1(
      dbg_0_dbg_uart_0_xfer_cnt[7]), .A2(dbg_0_dbg_uart_0_n_27_5));
  XNOR2_X1_LVT dbg_0_dbg_uart_0_i_27_15 (.ZN(dbg_0_dbg_uart_0_n_86), .A(
      dbg_0_dbg_uart_0_xfer_cnt[8]), .B(dbg_0_dbg_uart_0_n_27_6));
  NAND2_X1_LVT dbg_0_dbg_uart_0_i_31_26 (.ZN(dbg_0_dbg_uart_0_n_31_18), .A1(
      dbg_0_dbg_uart_0_n_96), .A2(dbg_0_dbg_uart_0_n_86));
  HA_X1_LVT dbg_0_dbg_uart_0_i_21_12 (.CO(dbg_0_dbg_uart_0_n_21_11), .S(
      dbg_0_dbg_uart_0_n_69), .A(dbg_0_dbg_uart_0_bit_cnt_max[9]), .B(
      dbg_0_dbg_uart_0_n_21_10));
  CLKGATETST_X1_LVT dbg_0_dbg_uart_0_clk_gate_sync_cnt_reg__5 (.GCK(
      dbg_0_dbg_uart_0_n_41), .CK(dbg_clk), .E(dbg_0_dbg_uart_0_n_76), .SE(1'b0));
  DFFS_X1_LVT \dbg_0_dbg_uart_0_sync_cnt_reg[12] (.Q(
      dbg_0_dbg_uart_0_bit_cnt_max[9]), .QN(), .CK(dbg_0_dbg_uart_0_n_41), .D(
      dbg_0_dbg_uart_0_n_69), .SN(dbg_0_dbg_uart_0_n_130));
  INV_X1_LVT dbg_0_dbg_uart_0_i_31_27 (.ZN(dbg_0_dbg_uart_0_n_31_19), .A(
      dbg_0_dbg_uart_0_bit_cnt_max[9]));
  OAI221_X1_LVT dbg_0_dbg_uart_0_i_31_28 (.ZN(dbg_0_dbg_uart_0_n_106), .A(
      dbg_0_dbg_uart_0_n_31_18), .B1(dbg_0_dbg_uart_0_n_31_2), .B2(
      dbg_0_dbg_uart_0_n_31_19), .C1(dbg_0_dbg_uart_0_n_31_5), .C2(
      dbg_0_dbg_uart_0_n_31_17));
  DFFR_X1_LVT \dbg_0_dbg_uart_0_xfer_cnt_reg[8] (.Q(dbg_0_dbg_uart_0_xfer_cnt[8]), 
      .QN(), .CK(dbg_0_dbg_uart_0_n_77), .D(dbg_0_dbg_uart_0_n_106), .RN(
      dbg_0_dbg_uart_0_n_130));
  OR2_X1_LVT dbg_0_dbg_uart_0_i_27_16 (.ZN(dbg_0_dbg_uart_0_n_27_7), .A1(
      dbg_0_dbg_uart_0_xfer_cnt[8]), .A2(dbg_0_dbg_uart_0_n_27_6));
  XNOR2_X1_LVT dbg_0_dbg_uart_0_i_27_17 (.ZN(dbg_0_dbg_uart_0_n_87), .A(
      dbg_0_dbg_uart_0_xfer_cnt[9]), .B(dbg_0_dbg_uart_0_n_27_7));
  NAND2_X1_LVT dbg_0_dbg_uart_0_i_31_29 (.ZN(dbg_0_dbg_uart_0_n_31_20), .A1(
      dbg_0_dbg_uart_0_n_96), .A2(dbg_0_dbg_uart_0_n_87));
  HA_X1_LVT dbg_0_dbg_uart_0_i_21_13 (.CO(dbg_0_dbg_uart_0_n_21_12), .S(
      dbg_0_dbg_uart_0_n_70), .A(dbg_0_dbg_uart_0_bit_cnt_max[10]), .B(
      dbg_0_dbg_uart_0_n_21_11));
  CLKGATETST_X1_LVT dbg_0_dbg_uart_0_clk_gate_sync_cnt_reg__4 (.GCK(
      dbg_0_dbg_uart_0_n_40), .CK(dbg_clk), .E(dbg_0_dbg_uart_0_n_76), .SE(1'b0));
  DFFS_X1_LVT \dbg_0_dbg_uart_0_sync_cnt_reg[13] (.Q(
      dbg_0_dbg_uart_0_bit_cnt_max[10]), .QN(), .CK(dbg_0_dbg_uart_0_n_40), .D(
      dbg_0_dbg_uart_0_n_70), .SN(dbg_0_dbg_uart_0_n_130));
  INV_X1_LVT dbg_0_dbg_uart_0_i_31_30 (.ZN(dbg_0_dbg_uart_0_n_31_21), .A(
      dbg_0_dbg_uart_0_bit_cnt_max[10]));
  OAI221_X1_LVT dbg_0_dbg_uart_0_i_31_31 (.ZN(dbg_0_dbg_uart_0_n_107), .A(
      dbg_0_dbg_uart_0_n_31_20), .B1(dbg_0_dbg_uart_0_n_31_2), .B2(
      dbg_0_dbg_uart_0_n_31_21), .C1(dbg_0_dbg_uart_0_n_31_5), .C2(
      dbg_0_dbg_uart_0_n_31_19));
  DFFR_X1_LVT \dbg_0_dbg_uart_0_xfer_cnt_reg[9] (.Q(dbg_0_dbg_uart_0_xfer_cnt[9]), 
      .QN(), .CK(dbg_0_dbg_uart_0_n_77), .D(dbg_0_dbg_uart_0_n_107), .RN(
      dbg_0_dbg_uart_0_n_130));
  OR2_X1_LVT dbg_0_dbg_uart_0_i_27_18 (.ZN(dbg_0_dbg_uart_0_n_27_8), .A1(
      dbg_0_dbg_uart_0_xfer_cnt[9]), .A2(dbg_0_dbg_uart_0_n_27_7));
  XNOR2_X1_LVT dbg_0_dbg_uart_0_i_27_19 (.ZN(dbg_0_dbg_uart_0_n_88), .A(
      dbg_0_dbg_uart_0_xfer_cnt[10]), .B(dbg_0_dbg_uart_0_n_27_8));
  NAND2_X1_LVT dbg_0_dbg_uart_0_i_31_32 (.ZN(dbg_0_dbg_uart_0_n_31_22), .A1(
      dbg_0_dbg_uart_0_n_96), .A2(dbg_0_dbg_uart_0_n_88));
  HA_X1_LVT dbg_0_dbg_uart_0_i_21_14 (.CO(dbg_0_dbg_uart_0_n_21_13), .S(
      dbg_0_dbg_uart_0_n_71), .A(dbg_0_dbg_uart_0_bit_cnt_max[11]), .B(
      dbg_0_dbg_uart_0_n_21_12));
  CLKGATETST_X1_LVT dbg_0_dbg_uart_0_clk_gate_sync_cnt_reg__3 (.GCK(
      dbg_0_dbg_uart_0_n_39), .CK(dbg_clk), .E(dbg_0_dbg_uart_0_n_76), .SE(1'b0));
  DFFS_X1_LVT \dbg_0_dbg_uart_0_sync_cnt_reg[14] (.Q(
      dbg_0_dbg_uart_0_bit_cnt_max[11]), .QN(), .CK(dbg_0_dbg_uart_0_n_39), .D(
      dbg_0_dbg_uart_0_n_71), .SN(dbg_0_dbg_uart_0_n_130));
  INV_X1_LVT dbg_0_dbg_uart_0_i_31_33 (.ZN(dbg_0_dbg_uart_0_n_31_23), .A(
      dbg_0_dbg_uart_0_bit_cnt_max[11]));
  OAI221_X1_LVT dbg_0_dbg_uart_0_i_31_34 (.ZN(dbg_0_dbg_uart_0_n_108), .A(
      dbg_0_dbg_uart_0_n_31_22), .B1(dbg_0_dbg_uart_0_n_31_2), .B2(
      dbg_0_dbg_uart_0_n_31_23), .C1(dbg_0_dbg_uart_0_n_31_5), .C2(
      dbg_0_dbg_uart_0_n_31_21));
  DFFR_X1_LVT \dbg_0_dbg_uart_0_xfer_cnt_reg[10] (.Q(
      dbg_0_dbg_uart_0_xfer_cnt[10]), .QN(), .CK(dbg_0_dbg_uart_0_n_77), .D(
      dbg_0_dbg_uart_0_n_108), .RN(dbg_0_dbg_uart_0_n_130));
  OR2_X1_LVT dbg_0_dbg_uart_0_i_27_20 (.ZN(dbg_0_dbg_uart_0_n_27_9), .A1(
      dbg_0_dbg_uart_0_xfer_cnt[10]), .A2(dbg_0_dbg_uart_0_n_27_8));
  XNOR2_X1_LVT dbg_0_dbg_uart_0_i_27_21 (.ZN(dbg_0_dbg_uart_0_n_89), .A(
      dbg_0_dbg_uart_0_xfer_cnt[11]), .B(dbg_0_dbg_uart_0_n_27_9));
  NAND2_X1_LVT dbg_0_dbg_uart_0_i_31_35 (.ZN(dbg_0_dbg_uart_0_n_31_24), .A1(
      dbg_0_dbg_uart_0_n_96), .A2(dbg_0_dbg_uart_0_n_89));
  HA_X1_LVT dbg_0_dbg_uart_0_i_21_15 (.CO(dbg_0_dbg_uart_0_n_21_14), .S(
      dbg_0_dbg_uart_0_n_72), .A(dbg_0_dbg_uart_0_bit_cnt_max[12]), .B(
      dbg_0_dbg_uart_0_n_21_13));
  CLKGATETST_X1_LVT dbg_0_dbg_uart_0_clk_gate_sync_cnt_reg__2 (.GCK(
      dbg_0_dbg_uart_0_n_38), .CK(dbg_clk), .E(dbg_0_dbg_uart_0_n_76), .SE(1'b0));
  DFFS_X1_LVT \dbg_0_dbg_uart_0_sync_cnt_reg[15] (.Q(
      dbg_0_dbg_uart_0_bit_cnt_max[12]), .QN(), .CK(dbg_0_dbg_uart_0_n_38), .D(
      dbg_0_dbg_uart_0_n_72), .SN(dbg_0_dbg_uart_0_n_130));
  INV_X1_LVT dbg_0_dbg_uart_0_i_31_36 (.ZN(dbg_0_dbg_uart_0_n_31_25), .A(
      dbg_0_dbg_uart_0_bit_cnt_max[12]));
  OAI221_X1_LVT dbg_0_dbg_uart_0_i_31_37 (.ZN(dbg_0_dbg_uart_0_n_109), .A(
      dbg_0_dbg_uart_0_n_31_24), .B1(dbg_0_dbg_uart_0_n_31_2), .B2(
      dbg_0_dbg_uart_0_n_31_25), .C1(dbg_0_dbg_uart_0_n_31_5), .C2(
      dbg_0_dbg_uart_0_n_31_23));
  DFFR_X1_LVT \dbg_0_dbg_uart_0_xfer_cnt_reg[11] (.Q(
      dbg_0_dbg_uart_0_xfer_cnt[11]), .QN(), .CK(dbg_0_dbg_uart_0_n_77), .D(
      dbg_0_dbg_uart_0_n_109), .RN(dbg_0_dbg_uart_0_n_130));
  NOR4_X1_LVT dbg_0_dbg_uart_0_i_32_2 (.ZN(dbg_0_dbg_uart_0_n_32_2), .A1(
      dbg_0_dbg_uart_0_xfer_cnt[8]), .A2(dbg_0_dbg_uart_0_xfer_cnt[9]), .A3(
      dbg_0_dbg_uart_0_xfer_cnt[10]), .A4(dbg_0_dbg_uart_0_xfer_cnt[11]));
  OR2_X1_LVT dbg_0_dbg_uart_0_i_27_22 (.ZN(dbg_0_dbg_uart_0_n_27_10), .A1(
      dbg_0_dbg_uart_0_xfer_cnt[11]), .A2(dbg_0_dbg_uart_0_n_27_9));
  XNOR2_X1_LVT dbg_0_dbg_uart_0_i_27_23 (.ZN(dbg_0_dbg_uart_0_n_90), .A(
      dbg_0_dbg_uart_0_xfer_cnt[12]), .B(dbg_0_dbg_uart_0_n_27_10));
  NAND2_X1_LVT dbg_0_dbg_uart_0_i_31_38 (.ZN(dbg_0_dbg_uart_0_n_31_26), .A1(
      dbg_0_dbg_uart_0_n_96), .A2(dbg_0_dbg_uart_0_n_90));
  HA_X1_LVT dbg_0_dbg_uart_0_i_21_16 (.CO(dbg_0_dbg_uart_0_n_21_15), .S(
      dbg_0_dbg_uart_0_n_73), .A(dbg_0_dbg_uart_0_bit_cnt_max[13]), .B(
      dbg_0_dbg_uart_0_n_21_14));
  CLKGATETST_X1_LVT dbg_0_dbg_uart_0_clk_gate_sync_cnt_reg__1 (.GCK(
      dbg_0_dbg_uart_0_n_37), .CK(dbg_clk), .E(dbg_0_dbg_uart_0_n_76), .SE(1'b0));
  DFFS_X1_LVT \dbg_0_dbg_uart_0_sync_cnt_reg[16] (.Q(
      dbg_0_dbg_uart_0_bit_cnt_max[13]), .QN(), .CK(dbg_0_dbg_uart_0_n_37), .D(
      dbg_0_dbg_uart_0_n_73), .SN(dbg_0_dbg_uart_0_n_130));
  INV_X1_LVT dbg_0_dbg_uart_0_i_31_39 (.ZN(dbg_0_dbg_uart_0_n_31_27), .A(
      dbg_0_dbg_uart_0_bit_cnt_max[13]));
  OAI221_X1_LVT dbg_0_dbg_uart_0_i_31_40 (.ZN(dbg_0_dbg_uart_0_n_110), .A(
      dbg_0_dbg_uart_0_n_31_26), .B1(dbg_0_dbg_uart_0_n_31_2), .B2(
      dbg_0_dbg_uart_0_n_31_27), .C1(dbg_0_dbg_uart_0_n_31_5), .C2(
      dbg_0_dbg_uart_0_n_31_25));
  DFFR_X1_LVT \dbg_0_dbg_uart_0_xfer_cnt_reg[12] (.Q(
      dbg_0_dbg_uart_0_xfer_cnt[12]), .QN(), .CK(dbg_0_dbg_uart_0_n_77), .D(
      dbg_0_dbg_uart_0_n_110), .RN(dbg_0_dbg_uart_0_n_130));
  OR2_X1_LVT dbg_0_dbg_uart_0_i_27_24 (.ZN(dbg_0_dbg_uart_0_n_27_11), .A1(
      dbg_0_dbg_uart_0_xfer_cnt[12]), .A2(dbg_0_dbg_uart_0_n_27_10));
  XNOR2_X1_LVT dbg_0_dbg_uart_0_i_27_25 (.ZN(dbg_0_dbg_uart_0_n_91), .A(
      dbg_0_dbg_uart_0_xfer_cnt[13]), .B(dbg_0_dbg_uart_0_n_27_11));
  NAND2_X1_LVT dbg_0_dbg_uart_0_i_31_41 (.ZN(dbg_0_dbg_uart_0_n_31_28), .A1(
      dbg_0_dbg_uart_0_n_96), .A2(dbg_0_dbg_uart_0_n_91));
  HA_X1_LVT dbg_0_dbg_uart_0_i_21_17 (.CO(dbg_0_dbg_uart_0_n_21_16), .S(
      dbg_0_dbg_uart_0_n_74), .A(dbg_0_dbg_uart_0_bit_cnt_max[14]), .B(
      dbg_0_dbg_uart_0_n_21_15));
  CLKGATETST_X1_LVT dbg_0_dbg_uart_0_clk_gate_sync_cnt_reg__0 (.GCK(
      dbg_0_dbg_uart_0_n_36), .CK(dbg_clk), .E(dbg_0_dbg_uart_0_n_76), .SE(1'b0));
  DFFS_X1_LVT \dbg_0_dbg_uart_0_sync_cnt_reg[17] (.Q(
      dbg_0_dbg_uart_0_bit_cnt_max[14]), .QN(), .CK(dbg_0_dbg_uart_0_n_36), .D(
      dbg_0_dbg_uart_0_n_74), .SN(dbg_0_dbg_uart_0_n_130));
  INV_X1_LVT dbg_0_dbg_uart_0_i_31_42 (.ZN(dbg_0_dbg_uart_0_n_31_29), .A(
      dbg_0_dbg_uart_0_bit_cnt_max[14]));
  OAI221_X1_LVT dbg_0_dbg_uart_0_i_31_43 (.ZN(dbg_0_dbg_uart_0_n_111), .A(
      dbg_0_dbg_uart_0_n_31_28), .B1(dbg_0_dbg_uart_0_n_31_2), .B2(
      dbg_0_dbg_uart_0_n_31_29), .C1(dbg_0_dbg_uart_0_n_31_5), .C2(
      dbg_0_dbg_uart_0_n_31_27));
  DFFR_X1_LVT \dbg_0_dbg_uart_0_xfer_cnt_reg[13] (.Q(
      dbg_0_dbg_uart_0_xfer_cnt[13]), .QN(), .CK(dbg_0_dbg_uart_0_n_77), .D(
      dbg_0_dbg_uart_0_n_111), .RN(dbg_0_dbg_uart_0_n_130));
  OR2_X1_LVT dbg_0_dbg_uart_0_i_27_26 (.ZN(dbg_0_dbg_uart_0_n_27_12), .A1(
      dbg_0_dbg_uart_0_xfer_cnt[13]), .A2(dbg_0_dbg_uart_0_n_27_11));
  XNOR2_X1_LVT dbg_0_dbg_uart_0_i_27_27 (.ZN(dbg_0_dbg_uart_0_n_92), .A(
      dbg_0_dbg_uart_0_xfer_cnt[14]), .B(dbg_0_dbg_uart_0_n_27_12));
  NAND2_X1_LVT dbg_0_dbg_uart_0_i_31_44 (.ZN(dbg_0_dbg_uart_0_n_31_30), .A1(
      dbg_0_dbg_uart_0_n_96), .A2(dbg_0_dbg_uart_0_n_92));
  XNOR2_X1_LVT dbg_0_dbg_uart_0_i_21_18 (.ZN(dbg_0_dbg_uart_0_n_21_17), .A(
      dbg_0_dbg_uart_0_bit_cnt_max[15]), .B(dbg_0_dbg_uart_0_n_21_16));
  INV_X1_LVT dbg_0_dbg_uart_0_i_21_19 (.ZN(dbg_0_dbg_uart_0_n_75), .A(
      dbg_0_dbg_uart_0_n_21_17));
  CLKGATETST_X1_LVT dbg_0_dbg_uart_0_clk_gate_sync_cnt_reg (.GCK(
      dbg_0_dbg_uart_0_n_35), .CK(dbg_clk), .E(dbg_0_dbg_uart_0_n_76), .SE(1'b0));
  DFFS_X1_LVT \dbg_0_dbg_uart_0_sync_cnt_reg[18] (.Q(
      dbg_0_dbg_uart_0_bit_cnt_max[15]), .QN(), .CK(dbg_0_dbg_uart_0_n_35), .D(
      dbg_0_dbg_uart_0_n_75), .SN(dbg_0_dbg_uart_0_n_130));
  INV_X1_LVT dbg_0_dbg_uart_0_i_31_45 (.ZN(dbg_0_dbg_uart_0_n_31_31), .A(
      dbg_0_dbg_uart_0_bit_cnt_max[15]));
  OAI221_X1_LVT dbg_0_dbg_uart_0_i_31_46 (.ZN(dbg_0_dbg_uart_0_n_112), .A(
      dbg_0_dbg_uart_0_n_31_30), .B1(dbg_0_dbg_uart_0_n_31_2), .B2(
      dbg_0_dbg_uart_0_n_31_31), .C1(dbg_0_dbg_uart_0_n_31_5), .C2(
      dbg_0_dbg_uart_0_n_31_29));
  DFFR_X1_LVT \dbg_0_dbg_uart_0_xfer_cnt_reg[14] (.Q(
      dbg_0_dbg_uart_0_xfer_cnt[14]), .QN(), .CK(dbg_0_dbg_uart_0_n_77), .D(
      dbg_0_dbg_uart_0_n_112), .RN(dbg_0_dbg_uart_0_n_130));
  OR2_X1_LVT dbg_0_dbg_uart_0_i_27_28 (.ZN(dbg_0_dbg_uart_0_n_27_13), .A1(
      dbg_0_dbg_uart_0_xfer_cnt[14]), .A2(dbg_0_dbg_uart_0_n_27_12));
  XNOR2_X1_LVT dbg_0_dbg_uart_0_i_27_29 (.ZN(dbg_0_dbg_uart_0_n_93), .A(
      dbg_0_dbg_uart_0_xfer_cnt[15]), .B(dbg_0_dbg_uart_0_n_27_13));
  AOI22_X1_LVT dbg_0_dbg_uart_0_i_31_47 (.ZN(dbg_0_dbg_uart_0_n_31_32), .A1(
      dbg_0_dbg_uart_0_n_97), .A2(dbg_0_dbg_uart_0_bit_cnt_max[15]), .B1(
      dbg_0_dbg_uart_0_n_96), .B2(dbg_0_dbg_uart_0_n_93));
  INV_X1_LVT dbg_0_dbg_uart_0_i_31_48 (.ZN(dbg_0_dbg_uart_0_n_113), .A(
      dbg_0_dbg_uart_0_n_31_32));
  DFFR_X1_LVT \dbg_0_dbg_uart_0_xfer_cnt_reg[15] (.Q(
      dbg_0_dbg_uart_0_xfer_cnt[15]), .QN(), .CK(dbg_0_dbg_uart_0_n_77), .D(
      dbg_0_dbg_uart_0_n_113), .RN(dbg_0_dbg_uart_0_n_130));
  NOR4_X1_LVT dbg_0_dbg_uart_0_i_32_3 (.ZN(dbg_0_dbg_uart_0_n_32_3), .A1(
      dbg_0_dbg_uart_0_xfer_cnt[12]), .A2(dbg_0_dbg_uart_0_xfer_cnt[13]), .A3(
      dbg_0_dbg_uart_0_xfer_cnt[14]), .A4(dbg_0_dbg_uart_0_xfer_cnt[15]));
  NAND4_X1_LVT dbg_0_dbg_uart_0_i_32_4 (.ZN(dbg_0_dbg_uart_0_n_114), .A1(
      dbg_0_dbg_uart_0_n_32_0), .A2(dbg_0_dbg_uart_0_n_32_1), .A3(
      dbg_0_dbg_uart_0_n_32_2), .A4(dbg_0_dbg_uart_0_n_32_3));
  NAND3_X1_LVT dbg_0_dbg_uart_0_i_33_2 (.ZN(dbg_0_dbg_uart_0_n_33_2), .A1(
      dbg_0_dbg_uart_0_n_33_0), .A2(dbg_0_dbg_uart_0_n_33_1), .A3(
      dbg_0_dbg_uart_0_n_114));
  NAND3_X1_LVT dbg_0_dbg_uart_0_i_33_3 (.ZN(dbg_0_dbg_uart_0_n_115), .A1(
      dbg_0_dbg_uart_0_n_33_2), .A2(dbg_0_dbg_uart_0_n_33_0), .A3(
      dbg_0_dbg_uart_0_n_33_1));
  CLKGATETST_X1_LVT dbg_0_dbg_uart_0_clk_gate_xfer_cnt_reg (.GCK(
      dbg_0_dbg_uart_0_n_77), .CK(dbg_clk), .E(dbg_0_dbg_uart_0_n_115), .SE(1'b0));
  DFFR_X1_LVT \dbg_0_dbg_uart_0_xfer_cnt_reg[0] (.Q(dbg_0_dbg_uart_0_xfer_cnt[0]), 
      .QN(), .CK(dbg_0_dbg_uart_0_n_77), .D(dbg_0_dbg_uart_0_n_98), .RN(
      dbg_0_dbg_uart_0_n_130));
  NOR4_X1_LVT dbg_0_dbg_uart_0_i_35_0 (.ZN(dbg_0_dbg_uart_0_n_35_0), .A1(
      dbg_0_dbg_uart_0_xfer_cnt[0]), .A2(dbg_0_dbg_uart_0_xfer_cnt[1]), .A3(
      dbg_0_dbg_uart_0_xfer_cnt[2]), .A4(dbg_0_dbg_uart_0_xfer_cnt[3]));
  NOR4_X1_LVT dbg_0_dbg_uart_0_i_35_1 (.ZN(dbg_0_dbg_uart_0_n_35_1), .A1(
      dbg_0_dbg_uart_0_xfer_cnt[4]), .A2(dbg_0_dbg_uart_0_xfer_cnt[5]), .A3(
      dbg_0_dbg_uart_0_xfer_cnt[6]), .A4(dbg_0_dbg_uart_0_xfer_cnt[7]));
  NOR4_X1_LVT dbg_0_dbg_uart_0_i_35_2 (.ZN(dbg_0_dbg_uart_0_n_35_2), .A1(
      dbg_0_dbg_uart_0_xfer_cnt[8]), .A2(dbg_0_dbg_uart_0_xfer_cnt[9]), .A3(
      dbg_0_dbg_uart_0_xfer_cnt[10]), .A4(dbg_0_dbg_uart_0_xfer_cnt[11]));
  NOR4_X1_LVT dbg_0_dbg_uart_0_i_35_3 (.ZN(dbg_0_dbg_uart_0_n_35_3), .A1(
      dbg_0_dbg_uart_0_xfer_cnt[12]), .A2(dbg_0_dbg_uart_0_xfer_cnt[13]), .A3(
      dbg_0_dbg_uart_0_xfer_cnt[14]), .A4(dbg_0_dbg_uart_0_xfer_cnt[15]));
  NAND4_X1_LVT dbg_0_dbg_uart_0_i_35_4 (.ZN(dbg_0_dbg_uart_0_n_35_4), .A1(
      dbg_0_dbg_uart_0_n_35_0), .A2(dbg_0_dbg_uart_0_n_35_1), .A3(
      dbg_0_dbg_uart_0_n_35_2), .A4(dbg_0_dbg_uart_0_n_35_3));
  NOR4_X1_LVT dbg_0_dbg_uart_0_i_35_5 (.ZN(dbg_0_dbg_uart_0_n_35_5), .A1(
      dbg_0_dbg_uart_0_xfer_bit[0]), .A2(dbg_0_dbg_uart_0_xfer_bit[1]), .A3(
      dbg_0_dbg_uart_0_xfer_bit[2]), .A4(dbg_0_dbg_uart_0_xfer_bit[3]));
  NOR2_X1_LVT dbg_0_dbg_uart_0_i_35_6 (.ZN(dbg_0_dbg_uart_0_xfer_bit_inc), .A1(
      dbg_0_dbg_uart_0_n_35_4), .A2(dbg_0_dbg_uart_0_n_35_5));
  INV_X1_LVT dbg_0_dbg_uart_0_i_5_1 (.ZN(dbg_0_dbg_uart_0_n_5_1), .A(
      dbg_0_dbg_uart_0_xfer_bit_inc));
  INV_X1_LVT dbg_0_dbg_uart_0_i_5_0 (.ZN(dbg_0_dbg_uart_0_n_5_0), .A(
      dbg_0_dbg_rd_rdy));
  NAND2_X1_LVT dbg_0_dbg_uart_0_i_5_2 (.ZN(dbg_0_dbg_uart_0_n_21), .A1(
      dbg_0_dbg_uart_0_n_5_1), .A2(dbg_0_dbg_uart_0_n_5_0));
  CLKGATETST_X1_LVT dbg_0_dbg_uart_0_clk_gate_xfer_buf_reg (.GCK(
      dbg_0_dbg_uart_0_n_0), .CK(dbg_clk), .E(dbg_0_dbg_uart_0_n_21), .SE(1'b0));
  DFFR_X1_LVT \dbg_0_dbg_uart_0_xfer_buf_reg[19] (.Q(
      dbg_0_dbg_uart_0_xfer_buf[19]), .QN(), .CK(dbg_0_dbg_uart_0_n_0), .D(
      dbg_0_dbg_uart_0_n_19), .RN(dbg_0_dbg_uart_0_n_130));
  AOI22_X1_LVT dbg_0_dbg_uart_0_i_4_34 (.ZN(dbg_0_dbg_uart_0_n_4_17), .A1(
      dbg_0_dbg_uart_0_n_4_0), .A2(dbg_0_dbg_uart_0_xfer_buf[19]), .B1(
      dbg_0_dbg_rd_rdy), .B2(dbg_0_dbg_dout[15]));
  INV_X1_LVT dbg_0_dbg_uart_0_i_4_35 (.ZN(dbg_0_dbg_uart_0_n_18), .A(
      dbg_0_dbg_uart_0_n_4_17));
  DFFR_X1_LVT \dbg_0_dbg_uart_0_xfer_buf_reg[18] (.Q(
      dbg_0_dbg_uart_0_xfer_buf[18]), .QN(), .CK(dbg_0_dbg_uart_0_n_0), .D(
      dbg_0_dbg_uart_0_n_18), .RN(dbg_0_dbg_uart_0_n_130));
  AOI22_X1_LVT dbg_0_dbg_uart_0_i_4_32 (.ZN(dbg_0_dbg_uart_0_n_4_16), .A1(
      dbg_0_dbg_uart_0_n_4_0), .A2(dbg_0_dbg_uart_0_xfer_buf[18]), .B1(
      dbg_0_dbg_rd_rdy), .B2(dbg_0_dbg_dout[14]));
  INV_X1_LVT dbg_0_dbg_uart_0_i_4_33 (.ZN(dbg_0_dbg_uart_0_n_17), .A(
      dbg_0_dbg_uart_0_n_4_16));
  DFFR_X1_LVT \dbg_0_dbg_uart_0_xfer_buf_reg[17] (.Q(
      dbg_0_dbg_uart_0_xfer_buf[17]), .QN(), .CK(dbg_0_dbg_uart_0_n_0), .D(
      dbg_0_dbg_uart_0_n_17), .RN(dbg_0_dbg_uart_0_n_130));
  AND2_X1_LVT dbg_0_dbg_uart_0_i_45_0 (.ZN(dbg_0_dbg_uart_0_cmd_valid), .A1(
      dbg_0_dbg_uart_0_n_27), .A2(dbg_0_dbg_uart_0_xfer_done));
  CLKGATETST_X1_LVT dbg_0_dbg_uart_0_clk_gate_dbg_addr_reg (.GCK(
      dbg_0_dbg_uart_0_n_129), .CK(dbg_clk), .E(dbg_0_dbg_uart_0_cmd_valid), .SE(
      1'b0));
  DFFR_X1_LVT \dbg_0_dbg_uart_0_dbg_addr_reg[5] (.Q(dbg_0_dbg_addr[5]), .QN(), 
      .CK(dbg_0_dbg_uart_0_n_129), .D(dbg_0_dbg_uart_0_xfer_buf[17]), .RN(
      dbg_0_dbg_uart_0_n_130));
  AOI22_X1_LVT dbg_0_dbg_uart_0_i_4_30 (.ZN(dbg_0_dbg_uart_0_n_4_15), .A1(
      dbg_0_dbg_uart_0_n_4_0), .A2(dbg_0_dbg_uart_0_xfer_buf[17]), .B1(
      dbg_0_dbg_rd_rdy), .B2(dbg_0_dbg_dout[13]));
  INV_X1_LVT dbg_0_dbg_uart_0_i_4_31 (.ZN(dbg_0_dbg_uart_0_n_16), .A(
      dbg_0_dbg_uart_0_n_4_15));
  DFFR_X1_LVT \dbg_0_dbg_uart_0_xfer_buf_reg[16] (.Q(
      dbg_0_dbg_uart_0_xfer_buf[16]), .QN(), .CK(dbg_0_dbg_uart_0_n_0), .D(
      dbg_0_dbg_uart_0_n_16), .RN(dbg_0_dbg_uart_0_n_130));
  DFFR_X1_LVT \dbg_0_dbg_uart_0_dbg_addr_reg[4] (.Q(dbg_0_dbg_addr[4]), .QN(), 
      .CK(dbg_0_dbg_uart_0_n_129), .D(dbg_0_dbg_uart_0_xfer_buf[16]), .RN(
      dbg_0_dbg_uart_0_n_130));
  AOI22_X1_LVT dbg_0_dbg_uart_0_i_4_28 (.ZN(dbg_0_dbg_uart_0_n_4_14), .A1(
      dbg_0_dbg_uart_0_n_4_0), .A2(dbg_0_dbg_uart_0_xfer_buf[16]), .B1(
      dbg_0_dbg_rd_rdy), .B2(dbg_0_dbg_dout[12]));
  INV_X1_LVT dbg_0_dbg_uart_0_i_4_29 (.ZN(dbg_0_dbg_uart_0_n_15), .A(
      dbg_0_dbg_uart_0_n_4_14));
  DFFR_X1_LVT \dbg_0_dbg_uart_0_xfer_buf_reg[15] (.Q(
      dbg_0_dbg_uart_0_xfer_buf[15]), .QN(), .CK(dbg_0_dbg_uart_0_n_0), .D(
      dbg_0_dbg_uart_0_n_15), .RN(dbg_0_dbg_uart_0_n_130));
  DFFR_X1_LVT \dbg_0_dbg_uart_0_dbg_addr_reg[3] (.Q(dbg_0_dbg_addr[3]), .QN(), 
      .CK(dbg_0_dbg_uart_0_n_129), .D(dbg_0_dbg_uart_0_xfer_buf[15]), .RN(
      dbg_0_dbg_uart_0_n_130));
  AOI22_X1_LVT dbg_0_dbg_uart_0_i_4_26 (.ZN(dbg_0_dbg_uart_0_n_4_13), .A1(
      dbg_0_dbg_uart_0_n_4_0), .A2(dbg_0_dbg_uart_0_xfer_buf[15]), .B1(
      dbg_0_dbg_rd_rdy), .B2(dbg_0_dbg_dout[11]));
  INV_X1_LVT dbg_0_dbg_uart_0_i_4_27 (.ZN(dbg_0_dbg_uart_0_n_14), .A(
      dbg_0_dbg_uart_0_n_4_13));
  DFFR_X1_LVT \dbg_0_dbg_uart_0_xfer_buf_reg[14] (.Q(
      dbg_0_dbg_uart_0_xfer_buf[14]), .QN(), .CK(dbg_0_dbg_uart_0_n_0), .D(
      dbg_0_dbg_uart_0_n_14), .RN(dbg_0_dbg_uart_0_n_130));
  DFFR_X1_LVT \dbg_0_dbg_uart_0_dbg_addr_reg[2] (.Q(dbg_0_dbg_addr[2]), .QN(), 
      .CK(dbg_0_dbg_uart_0_n_129), .D(dbg_0_dbg_uart_0_xfer_buf[14]), .RN(
      dbg_0_dbg_uart_0_n_130));
  AOI22_X1_LVT dbg_0_dbg_uart_0_i_4_24 (.ZN(dbg_0_dbg_uart_0_n_4_12), .A1(
      dbg_0_dbg_uart_0_n_4_0), .A2(dbg_0_dbg_uart_0_xfer_buf[14]), .B1(
      dbg_0_dbg_rd_rdy), .B2(dbg_0_dbg_dout[10]));
  INV_X1_LVT dbg_0_dbg_uart_0_i_4_25 (.ZN(dbg_0_dbg_uart_0_n_13), .A(
      dbg_0_dbg_uart_0_n_4_12));
  DFFR_X1_LVT \dbg_0_dbg_uart_0_xfer_buf_reg[13] (.Q(
      dbg_0_dbg_uart_0_xfer_buf[13]), .QN(), .CK(dbg_0_dbg_uart_0_n_0), .D(
      dbg_0_dbg_uart_0_n_13), .RN(dbg_0_dbg_uart_0_n_130));
  DFFR_X1_LVT \dbg_0_dbg_uart_0_dbg_addr_reg[1] (.Q(dbg_0_dbg_addr[1]), .QN(), 
      .CK(dbg_0_dbg_uart_0_n_129), .D(dbg_0_dbg_uart_0_xfer_buf[13]), .RN(
      dbg_0_dbg_uart_0_n_130));
  AOI22_X1_LVT dbg_0_dbg_uart_0_i_4_22 (.ZN(dbg_0_dbg_uart_0_n_4_11), .A1(
      dbg_0_dbg_uart_0_n_4_0), .A2(dbg_0_dbg_uart_0_xfer_buf[13]), .B1(
      dbg_0_dbg_rd_rdy), .B2(dbg_0_dbg_dout[9]));
  INV_X1_LVT dbg_0_dbg_uart_0_i_4_23 (.ZN(dbg_0_dbg_uart_0_n_12), .A(
      dbg_0_dbg_uart_0_n_4_11));
  DFFR_X1_LVT \dbg_0_dbg_uart_0_xfer_buf_reg[12] (.Q(
      dbg_0_dbg_uart_0_xfer_buf[12]), .QN(), .CK(dbg_0_dbg_uart_0_n_0), .D(
      dbg_0_dbg_uart_0_n_12), .RN(dbg_0_dbg_uart_0_n_130));
  DFFR_X1_LVT \dbg_0_dbg_uart_0_dbg_addr_reg[0] (.Q(dbg_0_dbg_addr[0]), .QN(), 
      .CK(dbg_0_dbg_uart_0_n_129), .D(dbg_0_dbg_uart_0_xfer_buf[12]), .RN(
      dbg_0_dbg_uart_0_n_130));
  INV_X1_LVT dbg_0_dbg_uart_0_i_49_0 (.ZN(dbg_0_dbg_uart_0_n_49_0), .A(
      dbg_0_mem_burst));
  CLKGATETST_X1_LVT dbg_0_dbg_uart_0_clk_gate_dbg_bw_reg (.GCK(
      dbg_0_dbg_uart_0_n_131), .CK(dbg_clk), .E(dbg_0_dbg_uart_0_cmd_valid), .SE(
      1'b0));
  DFFR_X1_LVT dbg_0_dbg_uart_0_dbg_bw_reg (.Q(dbg_0_dbg_uart_0_dbg_bw), .QN(), 
      .CK(dbg_0_dbg_uart_0_n_131), .D(dbg_0_dbg_uart_0_xfer_buf[18]), .RN(
      dbg_0_dbg_uart_0_n_130));
  AOI22_X1_LVT dbg_0_dbg_uart_0_i_49_1 (.ZN(dbg_0_dbg_uart_0_n_49_1), .A1(
      dbg_0_dbg_uart_0_n_49_0), .A2(dbg_0_dbg_uart_0_dbg_bw), .B1(
      dbg_0_mem_ctl[2]), .B2(dbg_0_mem_burst));
  AND2_X1_LVT dbg_0_dbg_uart_0_i_49_26 (.ZN(dbg_0_dbg_din[15]), .A1(
      dbg_0_dbg_uart_0_n_49_1), .A2(dbg_0_dbg_uart_0_xfer_buf[19]));
  AND2_X1_LVT dbg_0_dbg_uart_0_i_49_25 (.ZN(dbg_0_dbg_din[14]), .A1(
      dbg_0_dbg_uart_0_n_49_1), .A2(dbg_0_dbg_uart_0_xfer_buf[18]));
  AND2_X1_LVT dbg_0_dbg_uart_0_i_49_24 (.ZN(dbg_0_dbg_din[13]), .A1(
      dbg_0_dbg_uart_0_n_49_1), .A2(dbg_0_dbg_uart_0_xfer_buf[17]));
  AND2_X1_LVT dbg_0_dbg_uart_0_i_49_23 (.ZN(dbg_0_dbg_din[12]), .A1(
      dbg_0_dbg_uart_0_n_49_1), .A2(dbg_0_dbg_uart_0_xfer_buf[16]));
  AND2_X1_LVT dbg_0_dbg_uart_0_i_49_22 (.ZN(dbg_0_dbg_din[11]), .A1(
      dbg_0_dbg_uart_0_n_49_1), .A2(dbg_0_dbg_uart_0_xfer_buf[15]));
  AND2_X1_LVT dbg_0_dbg_uart_0_i_49_21 (.ZN(dbg_0_dbg_din[10]), .A1(
      dbg_0_dbg_uart_0_n_49_1), .A2(dbg_0_dbg_uart_0_xfer_buf[14]));
  AND2_X1_LVT dbg_0_dbg_uart_0_i_49_20 (.ZN(dbg_0_dbg_din[9]), .A1(
      dbg_0_dbg_uart_0_n_49_1), .A2(dbg_0_dbg_uart_0_xfer_buf[13]));
  AND2_X1_LVT dbg_0_dbg_uart_0_i_49_19 (.ZN(dbg_0_dbg_din[8]), .A1(
      dbg_0_dbg_uart_0_n_49_1), .A2(dbg_0_dbg_uart_0_xfer_buf[12]));
  INV_X1_LVT dbg_0_dbg_uart_0_i_49_2 (.ZN(dbg_0_dbg_uart_0_n_49_2), .A(
      dbg_0_dbg_uart_0_n_49_1));
  AOI22_X1_LVT dbg_0_dbg_uart_0_i_4_20 (.ZN(dbg_0_dbg_uart_0_n_4_10), .A1(
      dbg_0_dbg_uart_0_n_4_0), .A2(dbg_0_dbg_uart_0_xfer_buf[12]), .B1(
      dbg_0_dbg_rd_rdy), .B2(dbg_0_dbg_dout[8]));
  INV_X1_LVT dbg_0_dbg_uart_0_i_4_21 (.ZN(dbg_0_dbg_uart_0_n_11), .A(
      dbg_0_dbg_uart_0_n_4_10));
  DFFR_X1_LVT \dbg_0_dbg_uart_0_xfer_buf_reg[11] (.Q(
      dbg_0_dbg_uart_0_xfer_buf[11]), .QN(), .CK(dbg_0_dbg_uart_0_n_0), .D(
      dbg_0_dbg_uart_0_n_11), .RN(dbg_0_dbg_uart_0_n_130));
  AND2_X1_LVT dbg_0_dbg_uart_0_i_4_19 (.ZN(dbg_0_dbg_uart_0_n_10), .A1(
      dbg_0_dbg_uart_0_n_4_0), .A2(dbg_0_dbg_uart_0_xfer_buf[11]));
  DFFR_X1_LVT \dbg_0_dbg_uart_0_xfer_buf_reg[10] (.Q(
      dbg_0_dbg_uart_0_xfer_buf[10]), .QN(), .CK(dbg_0_dbg_uart_0_n_0), .D(
      dbg_0_dbg_uart_0_n_10), .RN(dbg_0_dbg_uart_0_n_130));
  AOI22_X1_LVT dbg_0_dbg_uart_0_i_49_17 (.ZN(dbg_0_dbg_uart_0_n_49_10), .A1(
      dbg_0_dbg_uart_0_n_49_2), .A2(dbg_0_dbg_uart_0_xfer_buf[19]), .B1(
      dbg_0_dbg_uart_0_n_49_1), .B2(dbg_0_dbg_uart_0_xfer_buf[10]));
  INV_X1_LVT dbg_0_dbg_uart_0_i_49_18 (.ZN(dbg_0_dbg_din[7]), .A(
      dbg_0_dbg_uart_0_n_49_10));
  INV_X1_LVT dbg_0_dbg_uart_0_i_4_18 (.ZN(dbg_0_dbg_uart_0_n_4_9), .A(
      dbg_0_dbg_uart_0_xfer_buf[10]));
  NAND2_X1_LVT dbg_0_dbg_uart_0_i_4_38 (.ZN(dbg_0_dbg_uart_0_n_20), .A1(
      dbg_0_dbg_uart_0_n_4_9), .A2(dbg_0_dbg_uart_0_n_4_0));
  DFFR_X1_LVT \dbg_0_dbg_uart_0_xfer_buf_reg[9] (.Q(dbg_0_dbg_uart_0_xfer_buf[9]), 
      .QN(), .CK(dbg_0_dbg_uart_0_n_0), .D(dbg_0_dbg_uart_0_n_20), .RN(
      dbg_0_dbg_uart_0_n_130));
  AOI22_X1_LVT dbg_0_dbg_uart_0_i_49_15 (.ZN(dbg_0_dbg_uart_0_n_49_9), .A1(
      dbg_0_dbg_uart_0_n_49_2), .A2(dbg_0_dbg_uart_0_xfer_buf[18]), .B1(
      dbg_0_dbg_uart_0_n_49_1), .B2(dbg_0_dbg_uart_0_xfer_buf[9]));
  INV_X1_LVT dbg_0_dbg_uart_0_i_49_16 (.ZN(dbg_0_dbg_din[6]), .A(
      dbg_0_dbg_uart_0_n_49_9));
  AOI22_X1_LVT dbg_0_dbg_uart_0_i_4_16 (.ZN(dbg_0_dbg_uart_0_n_4_8), .A1(
      dbg_0_dbg_uart_0_n_4_0), .A2(dbg_0_dbg_uart_0_xfer_buf[9]), .B1(
      dbg_0_dbg_rd_rdy), .B2(dbg_0_dbg_dout[7]));
  INV_X1_LVT dbg_0_dbg_uart_0_i_4_17 (.ZN(dbg_0_dbg_uart_0_n_9), .A(
      dbg_0_dbg_uart_0_n_4_8));
  DFFR_X1_LVT \dbg_0_dbg_uart_0_xfer_buf_reg[8] (.Q(dbg_0_dbg_uart_0_xfer_buf[8]), 
      .QN(), .CK(dbg_0_dbg_uart_0_n_0), .D(dbg_0_dbg_uart_0_n_9), .RN(
      dbg_0_dbg_uart_0_n_130));
  AOI22_X1_LVT dbg_0_dbg_uart_0_i_49_13 (.ZN(dbg_0_dbg_uart_0_n_49_8), .A1(
      dbg_0_dbg_uart_0_n_49_2), .A2(dbg_0_dbg_uart_0_xfer_buf[17]), .B1(
      dbg_0_dbg_uart_0_n_49_1), .B2(dbg_0_dbg_uart_0_xfer_buf[8]));
  INV_X1_LVT dbg_0_dbg_uart_0_i_49_14 (.ZN(dbg_0_dbg_din[5]), .A(
      dbg_0_dbg_uart_0_n_49_8));
  AOI22_X1_LVT dbg_0_dbg_uart_0_i_4_14 (.ZN(dbg_0_dbg_uart_0_n_4_7), .A1(
      dbg_0_dbg_uart_0_n_4_0), .A2(dbg_0_dbg_uart_0_xfer_buf[8]), .B1(
      dbg_0_dbg_rd_rdy), .B2(dbg_0_dbg_dout[6]));
  INV_X1_LVT dbg_0_dbg_uart_0_i_4_15 (.ZN(dbg_0_dbg_uart_0_n_8), .A(
      dbg_0_dbg_uart_0_n_4_7));
  DFFR_X1_LVT \dbg_0_dbg_uart_0_xfer_buf_reg[7] (.Q(dbg_0_dbg_uart_0_xfer_buf[7]), 
      .QN(), .CK(dbg_0_dbg_uart_0_n_0), .D(dbg_0_dbg_uart_0_n_8), .RN(
      dbg_0_dbg_uart_0_n_130));
  AOI22_X1_LVT dbg_0_dbg_uart_0_i_49_11 (.ZN(dbg_0_dbg_uart_0_n_49_7), .A1(
      dbg_0_dbg_uart_0_n_49_2), .A2(dbg_0_dbg_uart_0_xfer_buf[16]), .B1(
      dbg_0_dbg_uart_0_n_49_1), .B2(dbg_0_dbg_uart_0_xfer_buf[7]));
  INV_X1_LVT dbg_0_dbg_uart_0_i_49_12 (.ZN(dbg_0_dbg_din[4]), .A(
      dbg_0_dbg_uart_0_n_49_7));
  AOI22_X1_LVT dbg_0_dbg_uart_0_i_4_12 (.ZN(dbg_0_dbg_uart_0_n_4_6), .A1(
      dbg_0_dbg_uart_0_n_4_0), .A2(dbg_0_dbg_uart_0_xfer_buf[7]), .B1(
      dbg_0_dbg_rd_rdy), .B2(dbg_0_dbg_dout[5]));
  INV_X1_LVT dbg_0_dbg_uart_0_i_4_13 (.ZN(dbg_0_dbg_uart_0_n_7), .A(
      dbg_0_dbg_uart_0_n_4_6));
  DFFR_X1_LVT \dbg_0_dbg_uart_0_xfer_buf_reg[6] (.Q(dbg_0_dbg_uart_0_xfer_buf[6]), 
      .QN(), .CK(dbg_0_dbg_uart_0_n_0), .D(dbg_0_dbg_uart_0_n_7), .RN(
      dbg_0_dbg_uart_0_n_130));
  AOI22_X1_LVT dbg_0_dbg_uart_0_i_49_9 (.ZN(dbg_0_dbg_uart_0_n_49_6), .A1(
      dbg_0_dbg_uart_0_n_49_2), .A2(dbg_0_dbg_uart_0_xfer_buf[15]), .B1(
      dbg_0_dbg_uart_0_n_49_1), .B2(dbg_0_dbg_uart_0_xfer_buf[6]));
  INV_X1_LVT dbg_0_dbg_uart_0_i_49_10 (.ZN(dbg_0_dbg_din[3]), .A(
      dbg_0_dbg_uart_0_n_49_6));
  AOI22_X1_LVT dbg_0_dbg_uart_0_i_4_10 (.ZN(dbg_0_dbg_uart_0_n_4_5), .A1(
      dbg_0_dbg_uart_0_n_4_0), .A2(dbg_0_dbg_uart_0_xfer_buf[6]), .B1(
      dbg_0_dbg_rd_rdy), .B2(dbg_0_dbg_dout[4]));
  INV_X1_LVT dbg_0_dbg_uart_0_i_4_11 (.ZN(dbg_0_dbg_uart_0_n_6), .A(
      dbg_0_dbg_uart_0_n_4_5));
  DFFR_X1_LVT \dbg_0_dbg_uart_0_xfer_buf_reg[5] (.Q(dbg_0_dbg_uart_0_xfer_buf[5]), 
      .QN(), .CK(dbg_0_dbg_uart_0_n_0), .D(dbg_0_dbg_uart_0_n_6), .RN(
      dbg_0_dbg_uart_0_n_130));
  AOI22_X1_LVT dbg_0_dbg_uart_0_i_49_7 (.ZN(dbg_0_dbg_uart_0_n_49_5), .A1(
      dbg_0_dbg_uart_0_n_49_2), .A2(dbg_0_dbg_uart_0_xfer_buf[14]), .B1(
      dbg_0_dbg_uart_0_n_49_1), .B2(dbg_0_dbg_uart_0_xfer_buf[5]));
  INV_X1_LVT dbg_0_dbg_uart_0_i_49_8 (.ZN(dbg_0_dbg_din[2]), .A(
      dbg_0_dbg_uart_0_n_49_5));
  AOI22_X1_LVT dbg_0_dbg_uart_0_i_4_8 (.ZN(dbg_0_dbg_uart_0_n_4_4), .A1(
      dbg_0_dbg_uart_0_n_4_0), .A2(dbg_0_dbg_uart_0_xfer_buf[5]), .B1(
      dbg_0_dbg_rd_rdy), .B2(dbg_0_dbg_dout[3]));
  INV_X1_LVT dbg_0_dbg_uart_0_i_4_9 (.ZN(dbg_0_dbg_uart_0_n_5), .A(
      dbg_0_dbg_uart_0_n_4_4));
  DFFR_X1_LVT \dbg_0_dbg_uart_0_xfer_buf_reg[4] (.Q(dbg_0_dbg_uart_0_xfer_buf[4]), 
      .QN(), .CK(dbg_0_dbg_uart_0_n_0), .D(dbg_0_dbg_uart_0_n_5), .RN(
      dbg_0_dbg_uart_0_n_130));
  AOI22_X1_LVT dbg_0_dbg_uart_0_i_49_5 (.ZN(dbg_0_dbg_uart_0_n_49_4), .A1(
      dbg_0_dbg_uart_0_n_49_2), .A2(dbg_0_dbg_uart_0_xfer_buf[13]), .B1(
      dbg_0_dbg_uart_0_n_49_1), .B2(dbg_0_dbg_uart_0_xfer_buf[4]));
  INV_X1_LVT dbg_0_dbg_uart_0_i_49_6 (.ZN(dbg_0_dbg_din[1]), .A(
      dbg_0_dbg_uart_0_n_49_4));
  AOI22_X1_LVT dbg_0_dbg_uart_0_i_4_6 (.ZN(dbg_0_dbg_uart_0_n_4_3), .A1(
      dbg_0_dbg_uart_0_n_4_0), .A2(dbg_0_dbg_uart_0_xfer_buf[4]), .B1(
      dbg_0_dbg_rd_rdy), .B2(dbg_0_dbg_dout[2]));
  INV_X1_LVT dbg_0_dbg_uart_0_i_4_7 (.ZN(dbg_0_dbg_uart_0_n_4), .A(
      dbg_0_dbg_uart_0_n_4_3));
  DFFR_X1_LVT \dbg_0_dbg_uart_0_xfer_buf_reg[3] (.Q(dbg_0_dbg_uart_0_xfer_buf[3]), 
      .QN(), .CK(dbg_0_dbg_uart_0_n_0), .D(dbg_0_dbg_uart_0_n_4), .RN(
      dbg_0_dbg_uart_0_n_130));
  AOI22_X1_LVT dbg_0_dbg_uart_0_i_49_3 (.ZN(dbg_0_dbg_uart_0_n_49_3), .A1(
      dbg_0_dbg_uart_0_n_49_2), .A2(dbg_0_dbg_uart_0_xfer_buf[12]), .B1(
      dbg_0_dbg_uart_0_n_49_1), .B2(dbg_0_dbg_uart_0_xfer_buf[3]));
  INV_X1_LVT dbg_0_dbg_uart_0_i_49_4 (.ZN(dbg_0_dbg_din[0]), .A(
      dbg_0_dbg_uart_0_n_49_3));
  INV_X1_LVT dbg_0_dbg_uart_0_i_52_0 (.ZN(dbg_0_dbg_uart_0_n_52_0), .A(
      dbg_0_mem_burst));
  INV_X1_LVT dbg_0_dbg_uart_0_i_50_0 (.ZN(dbg_0_dbg_uart_0_n_50_0), .A(
      dbg_0_mem_burst_rd));
  INV_X1_LVT dbg_0_dbg_uart_0_i_50_1 (.ZN(dbg_0_dbg_uart_0_n_50_1), .A(
      dbg_0_dbg_uart_0_cmd_valid));
  OAI21_X1_LVT dbg_0_dbg_uart_0_i_50_2 (.ZN(dbg_0_dbg_uart_0_n_132), .A(
      dbg_0_dbg_uart_0_n_50_0), .B1(dbg_0_dbg_uart_0_n_50_1), .B2(
      dbg_0_dbg_uart_0_xfer_buf[19]));
  NOR3_X1_LVT dbg_0_dbg_uart_0_i_13_8 (.ZN(dbg_0_dbg_uart_0_n_30), .A1(
      dbg_0_dbg_uart_0_n_13_2), .A2(dbg_0_dbg_uart_0_n_13_1), .A3(
      dbg_0_dbg_uart_0_uart_state[1]));
  AND2_X1_LVT dbg_0_dbg_uart_0_i_51_0 (.ZN(dbg_0_dbg_uart_0_n_133), .A1(
      dbg_0_dbg_uart_0_xfer_done), .A2(dbg_0_dbg_uart_0_n_30));
  AOI22_X1_LVT dbg_0_dbg_uart_0_i_52_1 (.ZN(dbg_0_dbg_uart_0_n_52_1), .A1(
      dbg_0_dbg_uart_0_n_52_0), .A2(dbg_0_dbg_uart_0_n_132), .B1(
      dbg_0_dbg_uart_0_n_133), .B2(dbg_0_mem_burst));
  INV_X1_LVT dbg_0_dbg_uart_0_i_52_2 (.ZN(dbg_0_dbg_rd), .A(
      dbg_0_dbg_uart_0_n_52_1));
  AOI22_X1_LVT dbg_0_dbg_uart_0_i_4_4 (.ZN(dbg_0_dbg_uart_0_n_4_2), .A1(
      dbg_0_dbg_uart_0_n_4_0), .A2(dbg_0_dbg_uart_0_xfer_buf[3]), .B1(
      dbg_0_dbg_rd_rdy), .B2(dbg_0_dbg_dout[1]));
  INV_X1_LVT dbg_0_dbg_uart_0_i_4_5 (.ZN(dbg_0_dbg_uart_0_n_3), .A(
      dbg_0_dbg_uart_0_n_4_2));
  DFFR_X1_LVT \dbg_0_dbg_uart_0_xfer_buf_reg[2] (.Q(dbg_0_dbg_uart_0_xfer_buf[2]), 
      .QN(), .CK(dbg_0_dbg_uart_0_n_0), .D(dbg_0_dbg_uart_0_n_3), .RN(
      dbg_0_dbg_uart_0_n_130));
  AOI22_X1_LVT dbg_0_dbg_uart_0_i_4_2 (.ZN(dbg_0_dbg_uart_0_n_4_1), .A1(
      dbg_0_dbg_uart_0_n_4_0), .A2(dbg_0_dbg_uart_0_xfer_buf[2]), .B1(
      dbg_0_dbg_rd_rdy), .B2(dbg_0_dbg_dout[0]));
  INV_X1_LVT dbg_0_dbg_uart_0_i_4_3 (.ZN(dbg_0_dbg_uart_0_n_2), .A(
      dbg_0_dbg_uart_0_n_4_1));
  DFFR_X1_LVT \dbg_0_dbg_uart_0_xfer_buf_reg[1] (.Q(dbg_0_dbg_uart_0_xfer_buf[1]), 
      .QN(), .CK(dbg_0_dbg_uart_0_n_0), .D(dbg_0_dbg_uart_0_n_2), .RN(
      dbg_0_dbg_uart_0_n_130));
  AND2_X1_LVT dbg_0_dbg_uart_0_i_4_1 (.ZN(dbg_0_dbg_uart_0_n_1), .A1(
      dbg_0_dbg_uart_0_n_4_0), .A2(dbg_0_dbg_uart_0_xfer_buf[1]));
  DFFR_X1_LVT \dbg_0_dbg_uart_0_xfer_buf_reg[0] (.Q(dbg_0_dbg_uart_0_xfer_buf[0]), 
      .QN(), .CK(dbg_0_dbg_uart_0_n_0), .D(dbg_0_dbg_uart_0_n_1), .RN(
      dbg_0_dbg_uart_0_n_130));
  OAI21_X1_LVT dbg_0_dbg_uart_0_i_54_0 (.ZN(dbg_0_dbg_uart_0_n_54_0), .A(
      dbg_0_dbg_uart_0_xfer_bit_inc), .B1(dbg_0_dbg_uart_0_n_28), .B2(
      dbg_0_dbg_uart_0_n_30));
  INV_X1_LVT dbg_0_dbg_uart_0_i_54_1 (.ZN(dbg_0_dbg_uart_0_n_135), .A(
      dbg_0_dbg_uart_0_n_54_0));
  CLKGATETST_X1_LVT dbg_0_dbg_uart_0_clk_gate_dbg_uart_txd_reg (.GCK(
      dbg_0_dbg_uart_0_n_134), .CK(dbg_clk), .E(dbg_0_dbg_uart_0_n_135), .SE(
      1'b0));
  DFFS_X1_LVT dbg_0_dbg_uart_0_dbg_uart_txd_reg (.Q(dbg_uart_txd), .QN(), .CK(
      dbg_0_dbg_uart_0_n_134), .D(dbg_0_dbg_uart_0_xfer_buf[0]), .SN(
      dbg_0_dbg_uart_0_n_130));
  AND2_X1_LVT dbg_0_dbg_uart_0_i_56_0 (.ZN(dbg_0_dbg_wr), .A1(
      dbg_0_dbg_uart_0_xfer_done), .A2(dbg_0_dbg_uart_0_n_26));
  CLKGATETST_X1_LVT dbg_0_clk_gate_cpu_ctl_reg (.GCK(dbg_0_n_103), .CK(dbg_clk), 
      .E(dbg_0_cpu_ctl_wr), .SE(1'b0));
  DFFR_X1_LVT \dbg_0_cpu_ctl_reg[6] (.Q(dbg_cpu_reset), .QN(), .CK(dbg_0_n_103), 
      .D(dbg_0_dbg_din[6]), .RN(dbg_0_n_104));
  INV_X1_LVT dbg_0_i_53_0 (.ZN(dbg_0_n_53_0), .A(cpu_en_s));
  OAI21_X1_LVT dbg_0_i_53_1 (.ZN(dbg_0_n_53_1), .A(cpu_halt_st), .B1(
      dbg_0_n_53_0), .B2(dbg_0_cpu_ctl[1]));
  INV_X1_LVT dbg_0_i_53_2 (.ZN(dbg_freeze), .A(dbg_0_n_53_1));
  INV_X1_LVT dbg_0_i_55_0 (.ZN(dbg_0_n_55_0), .A(cpu_halt_st));
  NAND3_X1_LVT dbg_0_i_55_1 (.ZN(dbg_0_n_55_1), .A1(dbg_0_n_55_0), .A2(
      dbg_0_cpu_ctl_wr), .A3(dbg_0_dbg_din[0]));
  INV_X1_LVT dbg_0_i_55_2 (.ZN(dbg_0_n_55_2), .A(dbg_0_mem_state_nxt_reg[1]));
  NOR2_X1_LVT dbg_0_i_12_3 (.ZN(dbg_0_n_8), .A1(dbg_0_mem_state[0]), .A2(
      dbg_0_mem_state[1]));
  NAND3_X1_LVT dbg_0_i_55_3 (.ZN(dbg_0_n_55_3), .A1(dbg_0_n_55_2), .A2(
      dbg_0_mem_state_nxt_reg[0]), .A3(dbg_0_n_8));
  NAND3_X1_LVT dbg_0_i_55_4 (.ZN(dbg_0_n_55_4), .A1(puc_pnd_set), .A2(
      dbg_0_cpu_ctl[2]), .A3(dbg_en_s));
  INV_X1_LVT dbg_0_i_55_5 (.ZN(dbg_0_n_55_5), .A(dbg_0_dbg_swbrk));
  NAND4_X1_LVT dbg_0_i_55_6 (.ZN(dbg_0_halt_flag_set), .A1(dbg_0_n_55_1), .A2(
      dbg_0_n_55_3), .A3(dbg_0_n_55_4), .A4(dbg_0_n_55_5));
  INV_X1_LVT dbg_0_i_59_0 (.ZN(dbg_0_n_59_0), .A(dbg_0_halt_flag_set));
  INV_X1_LVT dbg_0_i_57_0 (.ZN(dbg_0_n_57_0), .A(dbg_0_n_7));
  NOR3_X1_LVT dbg_0_i_57_1 (.ZN(dbg_0_n_57_1), .A1(dbg_0_n_57_0), .A2(
      dbg_0_mem_state_nxt_reg[0]), .A3(dbg_0_mem_state_nxt_reg[1]));
  AND2_X1_LVT dbg_0_i_56_0 (.ZN(dbg_0_n_108), .A1(cpu_halt_st), .A2(
      dbg_0_cpu_ctl_wr));
  AOI21_X1_LVT dbg_0_i_57_2 (.ZN(dbg_0_n_57_2), .A(dbg_0_n_57_1), .B1(
      dbg_0_dbg_din[1]), .B2(dbg_0_n_108));
  INV_X1_LVT dbg_0_i_57_3 (.ZN(dbg_0_halt_flag_clr), .A(dbg_0_n_57_2));
  NOR2_X1_LVT dbg_0_i_59_1 (.ZN(dbg_0_n_110), .A1(dbg_0_n_59_0), .A2(
      dbg_0_halt_flag_clr));
  INV_X1_LVT dbg_0_i_60_1 (.ZN(dbg_0_n_60_1), .A(dbg_0_halt_flag_set));
  INV_X1_LVT dbg_0_i_60_0 (.ZN(dbg_0_n_60_0), .A(dbg_0_halt_flag_clr));
  NAND2_X1_LVT dbg_0_i_60_2 (.ZN(dbg_0_n_111), .A1(dbg_0_n_60_1), .A2(
      dbg_0_n_60_0));
  CLKGATETST_X1_LVT dbg_0_clk_gate_halt_flag_reg (.GCK(dbg_0_n_109), .CK(dbg_clk), 
      .E(dbg_0_n_111), .SE(1'b0));
  DFFR_X1_LVT dbg_0_halt_flag_reg (.Q(dbg_0_halt_flag), .QN(), .CK(dbg_0_n_109), 
      .D(dbg_0_n_110), .RN(dbg_0_n_104));
  NOR2_X1_LVT dbg_0_i_66_0 (.ZN(dbg_0_n_66_0), .A1(dbg_0_halt_flag), .A2(
      dbg_0_halt_flag_set));
  AND2_X1_LVT dbg_0_i_62_0 (.ZN(dbg_0_istep), .A1(dbg_0_dbg_din[2]), .A2(
      dbg_0_n_108));
  DFFR_X1_LVT \dbg_0_inc_step_reg[0] (.Q(dbg_0_n_113), .QN(), .CK(dbg_clk), .D(
      dbg_0_istep), .RN(dbg_0_n_104));
  INV_X1_LVT dbg_0_i_64_1 (.ZN(dbg_0_n_64_1), .A(dbg_0_n_113));
  INV_X1_LVT dbg_0_i_64_0 (.ZN(dbg_0_n_64_0), .A(dbg_0_istep));
  NAND2_X1_LVT dbg_0_i_64_2 (.ZN(dbg_0_n_114), .A1(dbg_0_n_64_1), .A2(
      dbg_0_n_64_0));
  DFFR_X1_LVT \dbg_0_inc_step_reg[1] (.Q(dbg_0_n_112), .QN(), .CK(dbg_clk), .D(
      dbg_0_n_114), .RN(dbg_0_n_104));
  NOR2_X1_LVT dbg_0_i_66_1 (.ZN(dbg_halt_cmd), .A1(dbg_0_n_66_0), .A2(
      dbg_0_n_112));
  NAND2_X1_LVT dbg_0_i_74_18 (.ZN(dbg_0_n_74_10), .A1(dbg_mem_addr[0]), .A2(
      dbg_0_mem_ctl[2]));
  INV_X1_LVT dbg_0_i_74_16 (.ZN(dbg_0_n_74_9), .A(dbg_0_mem_data[7]));
  INV_X1_LVT dbg_0_i_74_33 (.ZN(dbg_0_n_74_18), .A(dbg_0_mem_data[15]));
  OAI22_X1_LVT dbg_0_i_74_34 (.ZN(dbg_mem_dout[15]), .A1(dbg_0_n_74_10), .A2(
      dbg_0_n_74_9), .B1(dbg_0_mem_ctl[2]), .B2(dbg_0_n_74_18));
  INV_X1_LVT dbg_0_i_74_14 (.ZN(dbg_0_n_74_8), .A(dbg_0_mem_data[6]));
  INV_X1_LVT dbg_0_i_74_31 (.ZN(dbg_0_n_74_17), .A(dbg_0_mem_data[14]));
  OAI22_X1_LVT dbg_0_i_74_32 (.ZN(dbg_mem_dout[14]), .A1(dbg_0_n_74_10), .A2(
      dbg_0_n_74_8), .B1(dbg_0_mem_ctl[2]), .B2(dbg_0_n_74_17));
  INV_X1_LVT dbg_0_i_74_12 (.ZN(dbg_0_n_74_7), .A(dbg_0_mem_data[5]));
  INV_X1_LVT dbg_0_i_74_29 (.ZN(dbg_0_n_74_16), .A(dbg_0_mem_data[13]));
  OAI22_X1_LVT dbg_0_i_74_30 (.ZN(dbg_mem_dout[13]), .A1(dbg_0_n_74_10), .A2(
      dbg_0_n_74_7), .B1(dbg_0_mem_ctl[2]), .B2(dbg_0_n_74_16));
  INV_X1_LVT dbg_0_i_74_10 (.ZN(dbg_0_n_74_6), .A(dbg_0_mem_data[4]));
  INV_X1_LVT dbg_0_i_74_27 (.ZN(dbg_0_n_74_15), .A(dbg_0_mem_data[12]));
  OAI22_X1_LVT dbg_0_i_74_28 (.ZN(dbg_mem_dout[12]), .A1(dbg_0_n_74_10), .A2(
      dbg_0_n_74_6), .B1(dbg_0_mem_ctl[2]), .B2(dbg_0_n_74_15));
  INV_X1_LVT dbg_0_i_74_8 (.ZN(dbg_0_n_74_5), .A(dbg_0_mem_data[3]));
  INV_X1_LVT dbg_0_i_74_25 (.ZN(dbg_0_n_74_14), .A(dbg_0_mem_data[11]));
  OAI22_X1_LVT dbg_0_i_74_26 (.ZN(dbg_mem_dout[11]), .A1(dbg_0_n_74_10), .A2(
      dbg_0_n_74_5), .B1(dbg_0_mem_ctl[2]), .B2(dbg_0_n_74_14));
  INV_X1_LVT dbg_0_i_74_6 (.ZN(dbg_0_n_74_4), .A(dbg_0_mem_data[2]));
  INV_X1_LVT dbg_0_i_74_23 (.ZN(dbg_0_n_74_13), .A(dbg_0_mem_data[10]));
  OAI22_X1_LVT dbg_0_i_74_24 (.ZN(dbg_mem_dout[10]), .A1(dbg_0_n_74_10), .A2(
      dbg_0_n_74_4), .B1(dbg_0_mem_ctl[2]), .B2(dbg_0_n_74_13));
  INV_X1_LVT dbg_0_i_74_4 (.ZN(dbg_0_n_74_3), .A(dbg_0_mem_data[1]));
  INV_X1_LVT dbg_0_i_74_21 (.ZN(dbg_0_n_74_12), .A(dbg_0_mem_data[9]));
  OAI22_X1_LVT dbg_0_i_74_22 (.ZN(dbg_mem_dout[9]), .A1(dbg_0_n_74_10), .A2(
      dbg_0_n_74_3), .B1(dbg_0_mem_ctl[2]), .B2(dbg_0_n_74_12));
  INV_X1_LVT dbg_0_i_74_2 (.ZN(dbg_0_n_74_2), .A(dbg_0_mem_data[0]));
  INV_X1_LVT dbg_0_i_74_19 (.ZN(dbg_0_n_74_11), .A(dbg_0_mem_data[8]));
  OAI22_X1_LVT dbg_0_i_74_20 (.ZN(dbg_mem_dout[8]), .A1(dbg_0_n_74_10), .A2(
      dbg_0_n_74_2), .B1(dbg_0_mem_ctl[2]), .B2(dbg_0_n_74_11));
  INV_X1_LVT dbg_0_i_74_1 (.ZN(dbg_0_n_74_1), .A(dbg_mem_addr[0]));
  INV_X1_LVT dbg_0_i_74_0 (.ZN(dbg_0_n_74_0), .A(dbg_0_mem_ctl[2]));
  NOR2_X1_LVT dbg_0_i_74_35 (.ZN(dbg_0_n_74_19), .A1(dbg_0_n_74_1), .A2(
      dbg_0_n_74_0));
  NOR2_X1_LVT dbg_0_i_74_17 (.ZN(dbg_mem_dout[7]), .A1(dbg_0_n_74_19), .A2(
      dbg_0_n_74_9));
  NOR2_X1_LVT dbg_0_i_74_15 (.ZN(dbg_mem_dout[6]), .A1(dbg_0_n_74_19), .A2(
      dbg_0_n_74_8));
  NOR2_X1_LVT dbg_0_i_74_13 (.ZN(dbg_mem_dout[5]), .A1(dbg_0_n_74_19), .A2(
      dbg_0_n_74_7));
  NOR2_X1_LVT dbg_0_i_74_11 (.ZN(dbg_mem_dout[4]), .A1(dbg_0_n_74_19), .A2(
      dbg_0_n_74_6));
  NOR2_X1_LVT dbg_0_i_74_9 (.ZN(dbg_mem_dout[3]), .A1(dbg_0_n_74_19), .A2(
      dbg_0_n_74_5));
  NOR2_X1_LVT dbg_0_i_74_7 (.ZN(dbg_mem_dout[2]), .A1(dbg_0_n_74_19), .A2(
      dbg_0_n_74_4));
  NOR2_X1_LVT dbg_0_i_74_5 (.ZN(dbg_mem_dout[1]), .A1(dbg_0_n_74_19), .A2(
      dbg_0_n_74_3));
  NOR2_X1_LVT dbg_0_i_74_3 (.ZN(dbg_mem_dout[0]), .A1(dbg_0_n_74_19), .A2(
      dbg_0_n_74_2));
  OR2_X1_LVT multiplier_0_i_5_0 (.ZN(multiplier_0_n_15), .A1(per_we[0]), .A2(
      per_we[1]));
  NAND4_X1_LVT multiplier_0_i_0_0 (.ZN(multiplier_0_n_0_0), .A1(per_addr[3]), 
      .A2(per_addr[4]), .A3(per_addr[7]), .A4(per_en));
  NOR4_X1_LVT multiplier_0_i_0_1 (.ZN(multiplier_0_n_0_1), .A1(
      multiplier_0_n_0_0), .A2(per_addr[11]), .A3(per_addr[12]), .A4(
      per_addr[13]));
  NOR4_X1_LVT multiplier_0_i_0_2 (.ZN(multiplier_0_n_0_2), .A1(per_addr[6]), .A2(
      per_addr[8]), .A3(per_addr[9]), .A4(per_addr[10]));
  NAND2_X1_LVT multiplier_0_i_0_3 (.ZN(multiplier_0_n_0_3), .A1(
      multiplier_0_n_0_1), .A2(multiplier_0_n_0_2));
  NOR2_X1_LVT multiplier_0_i_0_4 (.ZN(multiplier_0_reg_sel), .A1(
      multiplier_0_n_0_3), .A2(per_addr[5]));
  AND2_X1_LVT multiplier_0_i_6_0 (.ZN(multiplier_0_reg_write), .A1(
      multiplier_0_n_15), .A2(multiplier_0_reg_sel));
  INV_X1_LVT multiplier_0_i_3_6 (.ZN(multiplier_0_n_3_2), .A(per_addr[2]));
  NOR3_X1_LVT multiplier_0_i_3_7 (.ZN(multiplier_0_n_5), .A1(multiplier_0_n_3_2), 
      .A2(per_addr[0]), .A3(per_addr[1]));
  AND2_X1_LVT multiplier_0_i_7_4 (.ZN(multiplier_0_op2_wr), .A1(
      multiplier_0_reg_write), .A2(multiplier_0_n_5));
  INV_X1_LVT multiplier_0_i_21_0 (.ZN(multiplier_0_n_38), .A(puc_rst));
  DFFR_X1_LVT \multiplier_0_cycle_reg[0] (.Q(multiplier_0_cycle[0]), .QN(), .CK(
      mclk), .D(multiplier_0_op2_wr), .RN(multiplier_0_n_38));
  DFFR_X1_LVT \multiplier_0_cycle_reg[1] (.Q(multiplier_0_cycle[1]), .QN(), .CK(
      mclk), .D(multiplier_0_cycle[0]), .RN(multiplier_0_n_38));
  INV_X1_LVT multiplier_0_i_60_0 (.ZN(multiplier_0_n_60_0), .A(
      multiplier_0_cycle[1]));
  INV_X1_LVT multiplier_0_i_38_0 (.ZN(multiplier_0_n_38_0), .A(
      multiplier_0_op2_wr));
  INV_X1_LVT multiplier_0_i_3_3 (.ZN(multiplier_0_n_3_1), .A(per_addr[1]));
  NOR3_X1_LVT multiplier_0_i_3_4 (.ZN(multiplier_0_n_3), .A1(multiplier_0_n_3_1), 
      .A2(per_addr[0]), .A3(per_addr[2]));
  AND2_X1_LVT multiplier_0_i_7_2 (.ZN(multiplier_0_n_18), .A1(
      multiplier_0_reg_write), .A2(multiplier_0_n_3));
  INV_X1_LVT multiplier_0_i_3_1 (.ZN(multiplier_0_n_3_0), .A(per_addr[0]));
  NOR3_X1_LVT multiplier_0_i_3_5 (.ZN(multiplier_0_n_4), .A1(multiplier_0_n_3_1), 
      .A2(multiplier_0_n_3_0), .A3(per_addr[2]));
  AND2_X1_LVT multiplier_0_i_7_3 (.ZN(multiplier_0_n_19), .A1(
      multiplier_0_reg_write), .A2(multiplier_0_n_4));
  OR2_X1_LVT multiplier_0_i_36_0 (.ZN(multiplier_0_n_68), .A1(multiplier_0_n_18), 
      .A2(multiplier_0_n_19));
  NOR3_X1_LVT multiplier_0_i_3_0 (.ZN(multiplier_0_n_1), .A1(per_addr[0]), .A2(
      per_addr[1]), .A3(per_addr[2]));
  AND2_X1_LVT multiplier_0_i_7_0 (.ZN(multiplier_0_n_16), .A1(multiplier_0_n_1), 
      .A2(multiplier_0_reg_write));
  NOR3_X1_LVT multiplier_0_i_3_2 (.ZN(multiplier_0_n_2), .A1(multiplier_0_n_3_0), 
      .A2(per_addr[1]), .A3(per_addr[2]));
  AND2_X1_LVT multiplier_0_i_7_1 (.ZN(multiplier_0_n_17), .A1(
      multiplier_0_reg_write), .A2(multiplier_0_n_2));
  OR4_X1_LVT multiplier_0_i_24_0 (.ZN(multiplier_0_op1_wr), .A1(
      multiplier_0_n_16), .A2(multiplier_0_n_19), .A3(multiplier_0_n_18), .A4(
      multiplier_0_n_17));
  CLKGATETST_X1_LVT multiplier_0_clk_gate_acc_sel_reg (.GCK(multiplier_0_n_67), 
      .CK(mclk), .E(multiplier_0_op1_wr), .SE(1'b0));
  DFFR_X1_LVT multiplier_0_acc_sel_reg (.Q(multiplier_0_acc_sel), .QN(), .CK(
      multiplier_0_n_67), .D(multiplier_0_n_68), .RN(multiplier_0_n_38));
  NOR2_X1_LVT multiplier_0_i_38_1 (.ZN(multiplier_0_result_clr), .A1(
      multiplier_0_n_38_0), .A2(multiplier_0_acc_sel));
  NOR3_X1_LVT multiplier_0_i_3_8 (.ZN(multiplier_0_n_6), .A1(multiplier_0_n_3_2), 
      .A2(multiplier_0_n_3_0), .A3(per_addr[1]));
  AND2_X1_LVT multiplier_0_i_7_5 (.ZN(multiplier_0_reslo_wr), .A1(
      multiplier_0_reg_write), .A2(multiplier_0_n_6));
  NOR2_X1_LVT multiplier_0_i_45_0 (.ZN(multiplier_0_n_45_0), .A1(
      multiplier_0_result_clr), .A2(multiplier_0_reslo_wr));
  INV_X1_LVT multiplier_0_i_34_16 (.ZN(multiplier_0_n_34_8), .A(
      multiplier_0_cycle[0]));
  INV_X1_LVT multiplier_0_i_29_0 (.ZN(multiplier_0_n_29_0), .A(
      multiplier_0_cycle[0]));
  CLKGATETST_X1_LVT multiplier_0_clk_gate_op2_reg (.GCK(multiplier_0_n_20), .CK(
      mclk), .E(multiplier_0_op2_wr), .SE(1'b0));
  DFFR_X1_LVT \multiplier_0_op2_reg[4] (.Q(multiplier_0_op2_reg[4]), .QN(), .CK(
      multiplier_0_n_20), .D(per_din[4]), .RN(multiplier_0_n_38));
  AND2_X1_LVT multiplier_0_i_8_4 (.ZN(multiplier_0_per_din_msk[12]), .A1(
      per_we[1]), .A2(per_din[12]));
  CLKGATETST_X1_LVT multiplier_0_clk_gate_op2_reg__0 (.GCK(multiplier_0_n_21), 
      .CK(mclk), .E(multiplier_0_op2_wr), .SE(1'b0));
  DFFR_X1_LVT \multiplier_0_op2_reg[12] (.Q(multiplier_0_op2_reg[12]), .QN(), 
      .CK(multiplier_0_n_21), .D(multiplier_0_per_din_msk[12]), .RN(
      multiplier_0_n_38));
  AOI22_X1_LVT multiplier_0_i_29_9 (.ZN(multiplier_0_n_29_5), .A1(
      multiplier_0_n_29_0), .A2(multiplier_0_op2_reg[4]), .B1(
      multiplier_0_cycle[0]), .B2(multiplier_0_op2_reg[12]));
  INV_X1_LVT multiplier_0_i_29_10 (.ZN(multiplier_0_op2_xp[4]), .A(
      multiplier_0_n_29_5));
  CLKGATETST_X1_LVT multiplier_0_clk_gate_op1_reg (.GCK(multiplier_0_n_41), .CK(
      mclk), .E(multiplier_0_op1_wr), .SE(1'b0));
  DFFR_X1_LVT \multiplier_0_op1_reg[3] (.Q(multiplier_0_op1[3]), .QN(), .CK(
      multiplier_0_n_41), .D(per_din[3]), .RN(multiplier_0_n_38));
  NAND2_X1_LVT multiplier_0_i_32_71 (.ZN(multiplier_0_n_32_71), .A1(
      multiplier_0_op2_xp[4]), .A2(multiplier_0_op1[3]));
  DFFR_X1_LVT \multiplier_0_op2_reg[3] (.Q(multiplier_0_op2_reg[3]), .QN(), .CK(
      multiplier_0_n_20), .D(per_din[3]), .RN(multiplier_0_n_38));
  AND2_X1_LVT multiplier_0_i_8_3 (.ZN(multiplier_0_per_din_msk[11]), .A1(
      per_we[1]), .A2(per_din[11]));
  DFFR_X1_LVT \multiplier_0_op2_reg[11] (.Q(multiplier_0_op2_reg[11]), .QN(), 
      .CK(multiplier_0_n_21), .D(multiplier_0_per_din_msk[11]), .RN(
      multiplier_0_n_38));
  AOI22_X1_LVT multiplier_0_i_29_7 (.ZN(multiplier_0_n_29_4), .A1(
      multiplier_0_n_29_0), .A2(multiplier_0_op2_reg[3]), .B1(
      multiplier_0_cycle[0]), .B2(multiplier_0_op2_reg[11]));
  INV_X1_LVT multiplier_0_i_29_8 (.ZN(multiplier_0_op2_xp[3]), .A(
      multiplier_0_n_29_4));
  DFFR_X1_LVT \multiplier_0_op1_reg[4] (.Q(multiplier_0_op1[4]), .QN(), .CK(
      multiplier_0_n_41), .D(per_din[4]), .RN(multiplier_0_n_38));
  NAND2_X1_LVT multiplier_0_i_32_55 (.ZN(multiplier_0_n_32_55), .A1(
      multiplier_0_op2_xp[3]), .A2(multiplier_0_op1[4]));
  XNOR2_X1_LVT multiplier_0_i_32_229 (.ZN(multiplier_0_n_32_234), .A(
      multiplier_0_n_32_71), .B(multiplier_0_n_32_55));
  DFFR_X1_LVT \multiplier_0_op2_reg[2] (.Q(multiplier_0_op2_reg[2]), .QN(), .CK(
      multiplier_0_n_20), .D(per_din[2]), .RN(multiplier_0_n_38));
  AND2_X1_LVT multiplier_0_i_8_2 (.ZN(multiplier_0_per_din_msk[10]), .A1(
      per_we[1]), .A2(per_din[10]));
  DFFR_X1_LVT \multiplier_0_op2_reg[10] (.Q(multiplier_0_op2_reg[10]), .QN(), 
      .CK(multiplier_0_n_21), .D(multiplier_0_per_din_msk[10]), .RN(
      multiplier_0_n_38));
  AOI22_X1_LVT multiplier_0_i_29_5 (.ZN(multiplier_0_n_29_3), .A1(
      multiplier_0_n_29_0), .A2(multiplier_0_op2_reg[2]), .B1(
      multiplier_0_cycle[0]), .B2(multiplier_0_op2_reg[10]));
  INV_X1_LVT multiplier_0_i_29_6 (.ZN(multiplier_0_op2_xp[2]), .A(
      multiplier_0_n_29_3));
  DFFR_X1_LVT \multiplier_0_op1_reg[5] (.Q(multiplier_0_op1[5]), .QN(), .CK(
      multiplier_0_n_41), .D(per_din[5]), .RN(multiplier_0_n_38));
  NAND2_X1_LVT multiplier_0_i_32_39 (.ZN(multiplier_0_n_32_39), .A1(
      multiplier_0_op2_xp[2]), .A2(multiplier_0_op1[5]));
  XNOR2_X1_LVT multiplier_0_i_32_230 (.ZN(multiplier_0_n_32_235), .A(
      multiplier_0_n_32_234), .B(multiplier_0_n_32_39));
  INV_X1_LVT multiplier_0_i_32_231 (.ZN(multiplier_0_n_32_236), .A(
      multiplier_0_n_32_235));
  DFFR_X1_LVT \multiplier_0_op2_reg[7] (.Q(multiplier_0_op2_reg[7]), .QN(), .CK(
      multiplier_0_n_20), .D(per_din[7]), .RN(multiplier_0_n_38));
  AND2_X1_LVT multiplier_0_i_8_7 (.ZN(multiplier_0_per_din_msk[15]), .A1(
      per_we[1]), .A2(per_din[15]));
  DFFR_X1_LVT \multiplier_0_op2_reg[15] (.Q(multiplier_0_op2_reg[15]), .QN(), 
      .CK(multiplier_0_n_21), .D(multiplier_0_per_din_msk[15]), .RN(
      multiplier_0_n_38));
  AOI22_X1_LVT multiplier_0_i_29_15 (.ZN(multiplier_0_n_29_8), .A1(
      multiplier_0_n_29_0), .A2(multiplier_0_op2_reg[7]), .B1(
      multiplier_0_cycle[0]), .B2(multiplier_0_op2_reg[15]));
  INV_X1_LVT multiplier_0_i_29_16 (.ZN(multiplier_0_op2_xp[7]), .A(
      multiplier_0_n_29_8));
  DFFR_X1_LVT \multiplier_0_op1_reg[0] (.Q(multiplier_0_op1[0]), .QN(), .CK(
      multiplier_0_n_41), .D(per_din[0]), .RN(multiplier_0_n_38));
  NAND2_X1_LVT multiplier_0_i_32_119 (.ZN(multiplier_0_n_32_119), .A1(
      multiplier_0_op2_xp[7]), .A2(multiplier_0_op1[0]));
  DFFR_X1_LVT \multiplier_0_op2_reg[6] (.Q(multiplier_0_op2_reg[6]), .QN(), .CK(
      multiplier_0_n_20), .D(per_din[6]), .RN(multiplier_0_n_38));
  AND2_X1_LVT multiplier_0_i_8_6 (.ZN(multiplier_0_per_din_msk[14]), .A1(
      per_we[1]), .A2(per_din[14]));
  DFFR_X1_LVT \multiplier_0_op2_reg[14] (.Q(multiplier_0_op2_reg[14]), .QN(), 
      .CK(multiplier_0_n_21), .D(multiplier_0_per_din_msk[14]), .RN(
      multiplier_0_n_38));
  AOI22_X1_LVT multiplier_0_i_29_13 (.ZN(multiplier_0_n_29_7), .A1(
      multiplier_0_n_29_0), .A2(multiplier_0_op2_reg[6]), .B1(
      multiplier_0_cycle[0]), .B2(multiplier_0_op2_reg[14]));
  INV_X1_LVT multiplier_0_i_29_14 (.ZN(multiplier_0_op2_xp[6]), .A(
      multiplier_0_n_29_7));
  DFFR_X1_LVT \multiplier_0_op1_reg[1] (.Q(multiplier_0_op1[1]), .QN(), .CK(
      multiplier_0_n_41), .D(per_din[1]), .RN(multiplier_0_n_38));
  NAND2_X1_LVT multiplier_0_i_32_103 (.ZN(multiplier_0_n_32_103), .A1(
      multiplier_0_op2_xp[6]), .A2(multiplier_0_op1[1]));
  XNOR2_X1_LVT multiplier_0_i_32_222 (.ZN(multiplier_0_n_32_227), .A(
      multiplier_0_n_32_119), .B(multiplier_0_n_32_103));
  DFFR_X1_LVT \multiplier_0_op2_reg[5] (.Q(multiplier_0_op2_reg[5]), .QN(), .CK(
      multiplier_0_n_20), .D(per_din[5]), .RN(multiplier_0_n_38));
  AND2_X1_LVT multiplier_0_i_8_5 (.ZN(multiplier_0_per_din_msk[13]), .A1(
      per_we[1]), .A2(per_din[13]));
  DFFR_X1_LVT \multiplier_0_op2_reg[13] (.Q(multiplier_0_op2_reg[13]), .QN(), 
      .CK(multiplier_0_n_21), .D(multiplier_0_per_din_msk[13]), .RN(
      multiplier_0_n_38));
  AOI22_X1_LVT multiplier_0_i_29_11 (.ZN(multiplier_0_n_29_6), .A1(
      multiplier_0_n_29_0), .A2(multiplier_0_op2_reg[5]), .B1(
      multiplier_0_cycle[0]), .B2(multiplier_0_op2_reg[13]));
  INV_X1_LVT multiplier_0_i_29_12 (.ZN(multiplier_0_op2_xp[5]), .A(
      multiplier_0_n_29_6));
  DFFR_X1_LVT \multiplier_0_op1_reg[2] (.Q(multiplier_0_op1[2]), .QN(), .CK(
      multiplier_0_n_41), .D(per_din[2]), .RN(multiplier_0_n_38));
  NAND2_X1_LVT multiplier_0_i_32_87 (.ZN(multiplier_0_n_32_87), .A1(
      multiplier_0_op2_xp[5]), .A2(multiplier_0_op1[2]));
  XNOR2_X1_LVT multiplier_0_i_32_223 (.ZN(multiplier_0_n_32_228), .A(
      multiplier_0_n_32_227), .B(multiplier_0_n_32_87));
  INV_X1_LVT multiplier_0_i_32_224 (.ZN(multiplier_0_n_32_229), .A(
      multiplier_0_n_32_228));
  NAND2_X1_LVT multiplier_0_i_32_85 (.ZN(multiplier_0_n_32_85), .A1(
      multiplier_0_op2_xp[5]), .A2(multiplier_0_op1[0]));
  NAND2_X1_LVT multiplier_0_i_32_69 (.ZN(multiplier_0_n_32_69), .A1(
      multiplier_0_op2_xp[4]), .A2(multiplier_0_op1[1]));
  XNOR2_X1_LVT multiplier_0_i_32_182 (.ZN(multiplier_0_n_32_183), .A(
      multiplier_0_n_32_85), .B(multiplier_0_n_32_69));
  NAND2_X1_LVT multiplier_0_i_32_53 (.ZN(multiplier_0_n_32_53), .A1(
      multiplier_0_op2_xp[3]), .A2(multiplier_0_op1[2]));
  XNOR2_X1_LVT multiplier_0_i_32_183 (.ZN(multiplier_0_n_32_184), .A(
      multiplier_0_n_32_183), .B(multiplier_0_n_32_53));
  INV_X1_LVT multiplier_0_i_32_184 (.ZN(multiplier_0_n_32_185), .A(
      multiplier_0_n_32_184));
  NAND2_X1_LVT multiplier_0_i_32_35 (.ZN(multiplier_0_n_32_35), .A1(
      multiplier_0_op2_xp[2]), .A2(multiplier_0_op1[1]));
  NAND2_X1_LVT multiplier_0_i_32_51 (.ZN(multiplier_0_n_32_51), .A1(
      multiplier_0_op2_xp[3]), .A2(multiplier_0_op1[0]));
  NOR2_X1_LVT multiplier_0_i_32_159 (.ZN(multiplier_0_n_32_159), .A1(
      multiplier_0_n_32_35), .A2(multiplier_0_n_32_51));
  DFFR_X1_LVT \multiplier_0_op2_reg[1] (.Q(multiplier_0_op2_reg[1]), .QN(), .CK(
      multiplier_0_n_20), .D(per_din[1]), .RN(multiplier_0_n_38));
  AND2_X1_LVT multiplier_0_i_8_1 (.ZN(multiplier_0_per_din_msk[9]), .A1(
      per_we[1]), .A2(per_din[9]));
  DFFR_X1_LVT \multiplier_0_op2_reg[9] (.Q(multiplier_0_op2_reg[9]), .QN(), .CK(
      multiplier_0_n_21), .D(multiplier_0_per_din_msk[9]), .RN(multiplier_0_n_38));
  AOI22_X1_LVT multiplier_0_i_29_3 (.ZN(multiplier_0_n_29_2), .A1(
      multiplier_0_n_29_0), .A2(multiplier_0_op2_reg[1]), .B1(
      multiplier_0_cycle[0]), .B2(multiplier_0_op2_reg[9]));
  INV_X1_LVT multiplier_0_i_29_4 (.ZN(multiplier_0_op2_xp[1]), .A(
      multiplier_0_n_29_2));
  NAND2_X1_LVT multiplier_0_i_32_19 (.ZN(multiplier_0_n_32_19), .A1(
      multiplier_0_op2_xp[1]), .A2(multiplier_0_op1[2]));
  NOR2_X1_LVT multiplier_0_i_32_160 (.ZN(multiplier_0_n_32_160), .A1(
      multiplier_0_n_32_19), .A2(multiplier_0_n_32_51));
  NOR2_X1_LVT multiplier_0_i_32_161 (.ZN(multiplier_0_n_32_161), .A1(
      multiplier_0_n_32_19), .A2(multiplier_0_n_32_35));
  OR3_X1_LVT multiplier_0_i_32_158 (.ZN(multiplier_0_n_32_158), .A1(
      multiplier_0_n_32_159), .A2(multiplier_0_n_32_160), .A3(
      multiplier_0_n_32_161));
  NAND2_X1_LVT multiplier_0_i_32_20 (.ZN(multiplier_0_n_32_20), .A1(
      multiplier_0_op2_xp[1]), .A2(multiplier_0_op1[3]));
  DFFR_X1_LVT \multiplier_0_op2_reg[0] (.Q(multiplier_0_op2_reg[0]), .QN(), .CK(
      multiplier_0_n_20), .D(per_din[0]), .RN(multiplier_0_n_38));
  AND2_X1_LVT multiplier_0_i_8_0 (.ZN(multiplier_0_per_din_msk[8]), .A1(
      per_din[8]), .A2(per_we[1]));
  DFFR_X1_LVT \multiplier_0_op2_reg[8] (.Q(multiplier_0_op2_reg[8]), .QN(), .CK(
      multiplier_0_n_21), .D(multiplier_0_per_din_msk[8]), .RN(multiplier_0_n_38));
  AOI22_X1_LVT multiplier_0_i_29_1 (.ZN(multiplier_0_n_29_1), .A1(
      multiplier_0_n_29_0), .A2(multiplier_0_op2_reg[0]), .B1(
      multiplier_0_op2_reg[8]), .B2(multiplier_0_cycle[0]));
  INV_X1_LVT multiplier_0_i_29_2 (.ZN(multiplier_0_op2_xp[0]), .A(
      multiplier_0_n_29_1));
  NAND2_X1_LVT multiplier_0_i_32_4 (.ZN(multiplier_0_n_32_4), .A1(
      multiplier_0_op2_xp[0]), .A2(multiplier_0_op1[4]));
  XNOR2_X1_LVT multiplier_0_i_32_173 (.ZN(multiplier_0_n_32_173), .A(
      multiplier_0_n_32_20), .B(multiplier_0_n_32_4));
  NAND2_X1_LVT multiplier_0_i_32_18 (.ZN(multiplier_0_n_32_18), .A1(
      multiplier_0_op2_xp[1]), .A2(multiplier_0_op1[1]));
  NAND2_X1_LVT multiplier_0_i_32_34 (.ZN(multiplier_0_n_32_34), .A1(
      multiplier_0_op2_xp[2]), .A2(multiplier_0_op1[0]));
  NOR2_X1_LVT multiplier_0_i_32_154 (.ZN(multiplier_0_n_32_154), .A1(
      multiplier_0_n_32_18), .A2(multiplier_0_n_32_34));
  NAND2_X1_LVT multiplier_0_i_32_3 (.ZN(multiplier_0_n_32_3), .A1(
      multiplier_0_op2_xp[0]), .A2(multiplier_0_op1[3]));
  INV_X1_LVT multiplier_0_i_32_164 (.ZN(multiplier_0_n_32_164), .A(
      multiplier_0_n_32_3));
  NAND2_X1_LVT multiplier_0_i_32_163 (.ZN(multiplier_0_n_32_163), .A1(
      multiplier_0_n_32_154), .A2(multiplier_0_n_32_164));
  INV_X1_LVT multiplier_0_i_32_165 (.ZN(multiplier_0_n_32_165), .A(
      multiplier_0_n_32_163));
  XNOR2_X1_LVT multiplier_0_i_32_174 (.ZN(multiplier_0_n_32_174), .A(
      multiplier_0_n_32_173), .B(multiplier_0_n_32_165));
  HA_X1_LVT multiplier_0_i_32_181 (.CO(multiplier_0_n_32_182), .S(
      multiplier_0_n_32_181), .A(multiplier_0_n_32_158), .B(
      multiplier_0_n_32_174));
  HA_X1_LVT multiplier_0_i_32_197 (.CO(multiplier_0_n_32_200), .S(
      multiplier_0_n_32_199), .A(multiplier_0_n_32_185), .B(
      multiplier_0_n_32_182));
  NAND2_X1_LVT multiplier_0_i_32_52 (.ZN(multiplier_0_n_32_52), .A1(
      multiplier_0_op2_xp[3]), .A2(multiplier_0_op1[1]));
  NAND2_X1_LVT multiplier_0_i_32_68 (.ZN(multiplier_0_n_32_68), .A1(
      multiplier_0_op2_xp[4]), .A2(multiplier_0_op1[0]));
  NOR2_X1_LVT multiplier_0_i_32_170 (.ZN(multiplier_0_n_32_170), .A1(
      multiplier_0_n_32_52), .A2(multiplier_0_n_32_68));
  NAND2_X1_LVT multiplier_0_i_32_36 (.ZN(multiplier_0_n_32_36), .A1(
      multiplier_0_op2_xp[2]), .A2(multiplier_0_op1[2]));
  NOR2_X1_LVT multiplier_0_i_32_171 (.ZN(multiplier_0_n_32_171), .A1(
      multiplier_0_n_32_36), .A2(multiplier_0_n_32_68));
  NOR2_X1_LVT multiplier_0_i_32_172 (.ZN(multiplier_0_n_32_172), .A1(
      multiplier_0_n_32_36), .A2(multiplier_0_n_32_52));
  OR3_X1_LVT multiplier_0_i_32_169 (.ZN(multiplier_0_n_32_169), .A1(
      multiplier_0_n_32_170), .A2(multiplier_0_n_32_171), .A3(
      multiplier_0_n_32_172));
  OR2_X1_LVT multiplier_0_i_32_176 (.ZN(multiplier_0_n_32_176), .A1(
      multiplier_0_n_32_4), .A2(multiplier_0_n_32_20));
  INV_X1_LVT multiplier_0_i_32_178 (.ZN(multiplier_0_n_32_178), .A(
      multiplier_0_n_32_20));
  NAND2_X1_LVT multiplier_0_i_32_177 (.ZN(multiplier_0_n_32_177), .A1(
      multiplier_0_n_32_165), .A2(multiplier_0_n_32_178));
  INV_X1_LVT multiplier_0_i_32_180 (.ZN(multiplier_0_n_32_180), .A(
      multiplier_0_n_32_4));
  NAND2_X1_LVT multiplier_0_i_32_179 (.ZN(multiplier_0_n_32_179), .A1(
      multiplier_0_n_32_165), .A2(multiplier_0_n_32_180));
  NAND3_X1_LVT multiplier_0_i_32_175 (.ZN(multiplier_0_n_32_175), .A1(
      multiplier_0_n_32_176), .A2(multiplier_0_n_32_177), .A3(
      multiplier_0_n_32_179));
  NAND2_X1_LVT multiplier_0_i_32_37 (.ZN(multiplier_0_n_32_37), .A1(
      multiplier_0_op2_xp[2]), .A2(multiplier_0_op1[3]));
  NAND2_X1_LVT multiplier_0_i_32_21 (.ZN(multiplier_0_n_32_21), .A1(
      multiplier_0_op2_xp[1]), .A2(multiplier_0_op1[4]));
  XNOR2_X1_LVT multiplier_0_i_32_189 (.ZN(multiplier_0_n_32_190), .A(
      multiplier_0_n_32_37), .B(multiplier_0_n_32_21));
  NAND2_X1_LVT multiplier_0_i_32_5 (.ZN(multiplier_0_n_32_5), .A1(
      multiplier_0_op2_xp[0]), .A2(multiplier_0_op1[5]));
  XNOR2_X1_LVT multiplier_0_i_32_190 (.ZN(multiplier_0_n_32_191), .A(
      multiplier_0_n_32_190), .B(multiplier_0_n_32_5));
  INV_X1_LVT multiplier_0_i_32_191 (.ZN(multiplier_0_n_32_192), .A(
      multiplier_0_n_32_191));
  FA_X1_LVT multiplier_0_i_32_196 (.CO(multiplier_0_n_32_198), .S(
      multiplier_0_n_32_197), .A(multiplier_0_n_32_169), .B(
      multiplier_0_n_32_175), .CI(multiplier_0_n_32_192));
  HA_X1_LVT multiplier_0_i_32_221 (.CO(multiplier_0_n_32_226), .S(
      multiplier_0_n_32_225), .A(multiplier_0_n_32_200), .B(
      multiplier_0_n_32_198));
  FA_X1_LVT multiplier_0_i_32_245 (.CO(multiplier_0_n_32_252), .S(
      multiplier_0_n_32_251), .A(multiplier_0_n_32_236), .B(
      multiplier_0_n_32_229), .CI(multiplier_0_n_32_226));
  NAND2_X1_LVT multiplier_0_i_32_86 (.ZN(multiplier_0_n_32_86), .A1(
      multiplier_0_op2_xp[5]), .A2(multiplier_0_op1[1]));
  NAND2_X1_LVT multiplier_0_i_32_102 (.ZN(multiplier_0_n_32_102), .A1(
      multiplier_0_op2_xp[6]), .A2(multiplier_0_op1[0]));
  NOR2_X1_LVT multiplier_0_i_32_202 (.ZN(multiplier_0_n_32_205), .A1(
      multiplier_0_n_32_86), .A2(multiplier_0_n_32_102));
  NAND2_X1_LVT multiplier_0_i_32_70 (.ZN(multiplier_0_n_32_70), .A1(
      multiplier_0_op2_xp[4]), .A2(multiplier_0_op1[2]));
  NOR2_X1_LVT multiplier_0_i_32_203 (.ZN(multiplier_0_n_32_206), .A1(
      multiplier_0_n_32_70), .A2(multiplier_0_n_32_102));
  NOR2_X1_LVT multiplier_0_i_32_204 (.ZN(multiplier_0_n_32_207), .A1(
      multiplier_0_n_32_70), .A2(multiplier_0_n_32_86));
  OR3_X1_LVT multiplier_0_i_32_201 (.ZN(multiplier_0_n_32_204), .A1(
      multiplier_0_n_32_205), .A2(multiplier_0_n_32_206), .A3(
      multiplier_0_n_32_207));
  NOR2_X1_LVT multiplier_0_i_32_193 (.ZN(multiplier_0_n_32_194), .A1(
      multiplier_0_n_32_21), .A2(multiplier_0_n_32_37));
  NOR2_X1_LVT multiplier_0_i_32_194 (.ZN(multiplier_0_n_32_195), .A1(
      multiplier_0_n_32_5), .A2(multiplier_0_n_32_37));
  NOR2_X1_LVT multiplier_0_i_32_195 (.ZN(multiplier_0_n_32_196), .A1(
      multiplier_0_n_32_5), .A2(multiplier_0_n_32_21));
  OR3_X1_LVT multiplier_0_i_32_192 (.ZN(multiplier_0_n_32_193), .A1(
      multiplier_0_n_32_194), .A2(multiplier_0_n_32_195), .A3(
      multiplier_0_n_32_196));
  DFFR_X1_LVT \multiplier_0_op1_reg[6] (.Q(multiplier_0_op1[6]), .QN(), .CK(
      multiplier_0_n_41), .D(per_din[6]), .RN(multiplier_0_n_38));
  NAND2_X1_LVT multiplier_0_i_32_6 (.ZN(multiplier_0_n_32_6), .A1(
      multiplier_0_op2_xp[0]), .A2(multiplier_0_op1[6]));
  INV_X1_LVT multiplier_0_i_32_217 (.ZN(multiplier_0_n_32_220), .A(
      multiplier_0_n_32_6));
  NAND2_X1_LVT multiplier_0_i_32_216 (.ZN(multiplier_0_n_32_219), .A1(
      multiplier_0_n_32_193), .A2(multiplier_0_n_32_220));
  NOR2_X1_LVT multiplier_0_i_32_186 (.ZN(multiplier_0_n_32_187), .A1(
      multiplier_0_n_32_69), .A2(multiplier_0_n_32_85));
  NOR2_X1_LVT multiplier_0_i_32_187 (.ZN(multiplier_0_n_32_188), .A1(
      multiplier_0_n_32_53), .A2(multiplier_0_n_32_85));
  NOR2_X1_LVT multiplier_0_i_32_188 (.ZN(multiplier_0_n_32_189), .A1(
      multiplier_0_n_32_53), .A2(multiplier_0_n_32_69));
  OR3_X1_LVT multiplier_0_i_32_185 (.ZN(multiplier_0_n_32_186), .A1(
      multiplier_0_n_32_187), .A2(multiplier_0_n_32_188), .A3(
      multiplier_0_n_32_189));
  NAND2_X1_LVT multiplier_0_i_32_218 (.ZN(multiplier_0_n_32_221), .A1(
      multiplier_0_n_32_186), .A2(multiplier_0_n_32_220));
  NAND2_X1_LVT multiplier_0_i_32_219 (.ZN(multiplier_0_n_32_222), .A1(
      multiplier_0_n_32_186), .A2(multiplier_0_n_32_193));
  NAND3_X1_LVT multiplier_0_i_32_215 (.ZN(multiplier_0_n_32_218), .A1(
      multiplier_0_n_32_219), .A2(multiplier_0_n_32_221), .A3(
      multiplier_0_n_32_222));
  NAND2_X1_LVT multiplier_0_i_32_23 (.ZN(multiplier_0_n_32_23), .A1(
      multiplier_0_op2_xp[1]), .A2(multiplier_0_op1[6]));
  DFFR_X1_LVT \multiplier_0_op1_reg[7] (.Q(multiplier_0_op1[7]), .QN(), .CK(
      multiplier_0_n_41), .D(per_din[7]), .RN(multiplier_0_n_38));
  NAND2_X1_LVT multiplier_0_i_32_7 (.ZN(multiplier_0_n_32_7), .A1(
      multiplier_0_op2_xp[0]), .A2(multiplier_0_op1[7]));
  XNOR2_X1_LVT multiplier_0_i_32_236 (.ZN(multiplier_0_n_32_241), .A(
      multiplier_0_n_32_23), .B(multiplier_0_n_32_7));
  NAND2_X1_LVT multiplier_0_i_32_38 (.ZN(multiplier_0_n_32_38), .A1(
      multiplier_0_op2_xp[2]), .A2(multiplier_0_op1[4]));
  NAND2_X1_LVT multiplier_0_i_32_54 (.ZN(multiplier_0_n_32_54), .A1(
      multiplier_0_op2_xp[3]), .A2(multiplier_0_op1[3]));
  NOR2_X1_LVT multiplier_0_i_32_209 (.ZN(multiplier_0_n_32_212), .A1(
      multiplier_0_n_32_38), .A2(multiplier_0_n_32_54));
  NAND2_X1_LVT multiplier_0_i_32_22 (.ZN(multiplier_0_n_32_22), .A1(
      multiplier_0_op2_xp[1]), .A2(multiplier_0_op1[5]));
  NOR2_X1_LVT multiplier_0_i_32_210 (.ZN(multiplier_0_n_32_213), .A1(
      multiplier_0_n_32_22), .A2(multiplier_0_n_32_54));
  NOR2_X1_LVT multiplier_0_i_32_211 (.ZN(multiplier_0_n_32_214), .A1(
      multiplier_0_n_32_22), .A2(multiplier_0_n_32_38));
  OR3_X1_LVT multiplier_0_i_32_208 (.ZN(multiplier_0_n_32_211), .A1(
      multiplier_0_n_32_212), .A2(multiplier_0_n_32_213), .A3(
      multiplier_0_n_32_214));
  XNOR2_X1_LVT multiplier_0_i_32_237 (.ZN(multiplier_0_n_32_242), .A(
      multiplier_0_n_32_241), .B(multiplier_0_n_32_211));
  FA_X1_LVT multiplier_0_i_32_244 (.CO(multiplier_0_n_32_250), .S(
      multiplier_0_n_32_249), .A(multiplier_0_n_32_204), .B(
      multiplier_0_n_32_218), .CI(multiplier_0_n_32_242));
  XNOR2_X1_LVT multiplier_0_i_32_205 (.ZN(multiplier_0_n_32_208), .A(
      multiplier_0_n_32_54), .B(multiplier_0_n_32_38));
  XNOR2_X1_LVT multiplier_0_i_32_206 (.ZN(multiplier_0_n_32_209), .A(
      multiplier_0_n_32_208), .B(multiplier_0_n_32_22));
  INV_X1_LVT multiplier_0_i_32_207 (.ZN(multiplier_0_n_32_210), .A(
      multiplier_0_n_32_209));
  XNOR2_X1_LVT multiplier_0_i_32_198 (.ZN(multiplier_0_n_32_201), .A(
      multiplier_0_n_32_102), .B(multiplier_0_n_32_86));
  XNOR2_X1_LVT multiplier_0_i_32_199 (.ZN(multiplier_0_n_32_202), .A(
      multiplier_0_n_32_201), .B(multiplier_0_n_32_70));
  INV_X1_LVT multiplier_0_i_32_200 (.ZN(multiplier_0_n_32_203), .A(
      multiplier_0_n_32_202));
  XNOR2_X1_LVT multiplier_0_i_32_212 (.ZN(multiplier_0_n_32_215), .A(
      multiplier_0_n_32_6), .B(multiplier_0_n_32_193));
  XNOR2_X1_LVT multiplier_0_i_32_213 (.ZN(multiplier_0_n_32_216), .A(
      multiplier_0_n_32_215), .B(multiplier_0_n_32_186));
  INV_X1_LVT multiplier_0_i_32_214 (.ZN(multiplier_0_n_32_217), .A(
      multiplier_0_n_32_216));
  FA_X1_LVT multiplier_0_i_32_220 (.CO(multiplier_0_n_32_224), .S(
      multiplier_0_n_32_223), .A(multiplier_0_n_32_210), .B(
      multiplier_0_n_32_203), .CI(multiplier_0_n_32_217));
  HA_X1_LVT multiplier_0_i_32_246 (.CO(multiplier_0_n_32_254), .S(
      multiplier_0_n_32_253), .A(multiplier_0_n_32_249), .B(
      multiplier_0_n_32_224));
  XNOR2_X1_LVT multiplier_0_i_32_166 (.ZN(multiplier_0_n_32_166), .A(
      multiplier_0_n_32_68), .B(multiplier_0_n_32_52));
  XNOR2_X1_LVT multiplier_0_i_32_167 (.ZN(multiplier_0_n_32_167), .A(
      multiplier_0_n_32_166), .B(multiplier_0_n_32_36));
  INV_X1_LVT multiplier_0_i_32_168 (.ZN(multiplier_0_n_32_168), .A(
      multiplier_0_n_32_167));
  XNOR2_X1_LVT multiplier_0_i_32_162 (.ZN(multiplier_0_n_32_162), .A(
      multiplier_0_n_32_3), .B(multiplier_0_n_32_154));
  XNOR2_X1_LVT multiplier_0_i_32_155 (.ZN(multiplier_0_n_32_155), .A(
      multiplier_0_n_32_51), .B(multiplier_0_n_32_35));
  XNOR2_X1_LVT multiplier_0_i_32_156 (.ZN(multiplier_0_n_32_156), .A(
      multiplier_0_n_32_155), .B(multiplier_0_n_32_19));
  INV_X1_LVT multiplier_0_i_32_157 (.ZN(multiplier_0_n_32_157), .A(
      multiplier_0_n_32_156));
  XNOR2_X1_LVT multiplier_0_i_32_152 (.ZN(multiplier_0_n_32_152), .A(
      multiplier_0_n_32_34), .B(multiplier_0_n_32_18));
  INV_X1_LVT multiplier_0_i_32_153 (.ZN(multiplier_0_n_32_153), .A(
      multiplier_0_n_32_152));
  NAND2_X1_LVT multiplier_0_i_32_2 (.ZN(multiplier_0_n_32_2), .A1(
      multiplier_0_op2_xp[0]), .A2(multiplier_0_op1[2]));
  INV_X1_LVT multiplier_0_i_32_594 (.ZN(multiplier_0_n_32_651), .A(
      multiplier_0_n_32_2));
  NAND2_X1_LVT multiplier_0_i_32_593 (.ZN(multiplier_0_n_32_650), .A1(
      multiplier_0_n_32_153), .A2(multiplier_0_n_32_651));
  NAND2_X1_LVT multiplier_0_i_32_1 (.ZN(multiplier_0_n_32_1), .A1(
      multiplier_0_op2_xp[0]), .A2(multiplier_0_op1[1]));
  NAND2_X1_LVT multiplier_0_i_32_17 (.ZN(multiplier_0_n_32_17), .A1(
      multiplier_0_op2_xp[1]), .A2(multiplier_0_op1[0]));
  NOR2_X1_LVT multiplier_0_i_32_588 (.ZN(multiplier_0_n_32_646), .A1(
      multiplier_0_n_32_1), .A2(multiplier_0_n_32_17));
  NAND2_X1_LVT multiplier_0_i_32_595 (.ZN(multiplier_0_n_32_652), .A1(
      multiplier_0_n_32_646), .A2(multiplier_0_n_32_651));
  NAND2_X1_LVT multiplier_0_i_32_596 (.ZN(multiplier_0_n_32_653), .A1(
      multiplier_0_n_32_646), .A2(multiplier_0_n_32_153));
  NAND3_X1_LVT multiplier_0_i_32_592 (.ZN(multiplier_0_n_32_649), .A1(
      multiplier_0_n_32_650), .A2(multiplier_0_n_32_652), .A3(
      multiplier_0_n_32_653));
  FA_X1_LVT multiplier_0_i_32_597 (.CO(multiplier_0_n_32_654), .S(
      multiplier_0_n_45), .A(multiplier_0_n_32_162), .B(multiplier_0_n_32_157), 
      .CI(multiplier_0_n_32_649));
  FA_X1_LVT multiplier_0_i_32_598 (.CO(multiplier_0_n_32_655), .S(
      multiplier_0_n_46), .A(multiplier_0_n_32_168), .B(multiplier_0_n_32_181), 
      .CI(multiplier_0_n_32_654));
  FA_X1_LVT multiplier_0_i_32_599 (.CO(multiplier_0_n_32_656), .S(
      multiplier_0_n_47), .A(multiplier_0_n_32_197), .B(multiplier_0_n_32_199), 
      .CI(multiplier_0_n_32_655));
  FA_X1_LVT multiplier_0_i_32_600 (.CO(multiplier_0_n_32_657), .S(
      multiplier_0_n_48), .A(multiplier_0_n_32_225), .B(multiplier_0_n_32_223), 
      .CI(multiplier_0_n_32_656));
  FA_X1_LVT multiplier_0_i_32_601 (.CO(multiplier_0_n_32_658), .S(
      multiplier_0_n_49), .A(multiplier_0_n_32_251), .B(multiplier_0_n_32_253), 
      .CI(multiplier_0_n_32_657));
  INV_X1_LVT multiplier_0_i_34_14 (.ZN(multiplier_0_n_34_7), .A(
      multiplier_0_n_49));
  OR2_X1_LVT multiplier_0_i_26_0 (.ZN(multiplier_0_n_40), .A1(multiplier_0_n_17), 
      .A2(multiplier_0_n_19));
  CLKGATETST_X1_LVT multiplier_0_clk_gate_sign_sel_reg (.GCK(multiplier_0_n_39), 
      .CK(mclk), .E(multiplier_0_op1_wr), .SE(1'b0));
  DFFR_X1_LVT multiplier_0_sign_sel_reg (.Q(multiplier_0_sign_sel), .QN(), .CK(
      multiplier_0_n_39), .D(multiplier_0_n_40), .RN(multiplier_0_n_38));
  AND2_X1_LVT multiplier_0_i_28_0 (.ZN(multiplier_0_op2_hi_xp[8]), .A1(
      multiplier_0_op2_reg[15]), .A2(multiplier_0_sign_sel));
  AND2_X1_LVT multiplier_0_i_29_17 (.ZN(multiplier_0_op2_xp[8]), .A1(
      multiplier_0_cycle[0]), .A2(multiplier_0_op2_hi_xp[8]));
  NAND2_X1_LVT multiplier_0_i_32_141 (.ZN(multiplier_0_n_32_141), .A1(
      multiplier_0_op2_xp[8]), .A2(multiplier_0_op1[5]));
  NAND2_X1_LVT multiplier_0_i_32_125 (.ZN(multiplier_0_n_32_125), .A1(
      multiplier_0_op2_xp[7]), .A2(multiplier_0_op1[6]));
  XNOR2_X1_LVT multiplier_0_i_32_380 (.ZN(multiplier_0_n_32_407), .A(
      multiplier_0_n_32_141), .B(multiplier_0_n_32_125));
  NAND2_X1_LVT multiplier_0_i_32_109 (.ZN(multiplier_0_n_32_109), .A1(
      multiplier_0_op2_xp[6]), .A2(multiplier_0_op1[7]));
  XNOR2_X1_LVT multiplier_0_i_32_381 (.ZN(multiplier_0_n_32_408), .A(
      multiplier_0_n_32_407), .B(multiplier_0_n_32_109));
  DFFR_X1_LVT \multiplier_0_op1_reg[11] (.Q(multiplier_0_op1[11]), .QN(), .CK(
      multiplier_0_n_41), .D(multiplier_0_per_din_msk[11]), .RN(
      multiplier_0_n_38));
  NAND2_X1_LVT multiplier_0_i_32_28 (.ZN(multiplier_0_n_32_28), .A1(
      multiplier_0_op2_xp[1]), .A2(multiplier_0_op1[11]));
  DFFR_X1_LVT \multiplier_0_op1_reg[10] (.Q(multiplier_0_op1[10]), .QN(), .CK(
      multiplier_0_n_41), .D(multiplier_0_per_din_msk[10]), .RN(
      multiplier_0_n_38));
  NAND2_X1_LVT multiplier_0_i_32_44 (.ZN(multiplier_0_n_32_44), .A1(
      multiplier_0_op2_xp[2]), .A2(multiplier_0_op1[10]));
  NOR2_X1_LVT multiplier_0_i_32_373 (.ZN(multiplier_0_n_32_396), .A1(
      multiplier_0_n_32_28), .A2(multiplier_0_n_32_44));
  DFFR_X1_LVT \multiplier_0_op1_reg[12] (.Q(multiplier_0_op1[12]), .QN(), .CK(
      multiplier_0_n_41), .D(multiplier_0_per_din_msk[12]), .RN(
      multiplier_0_n_38));
  NAND2_X1_LVT multiplier_0_i_32_12 (.ZN(multiplier_0_n_32_12), .A1(
      multiplier_0_op2_xp[0]), .A2(multiplier_0_op1[12]));
  NOR2_X1_LVT multiplier_0_i_32_374 (.ZN(multiplier_0_n_32_397), .A1(
      multiplier_0_n_32_12), .A2(multiplier_0_n_32_44));
  NOR2_X1_LVT multiplier_0_i_32_375 (.ZN(multiplier_0_n_32_398), .A1(
      multiplier_0_n_32_12), .A2(multiplier_0_n_32_28));
  OR3_X1_LVT multiplier_0_i_32_372 (.ZN(multiplier_0_n_32_395), .A1(
      multiplier_0_n_32_396), .A2(multiplier_0_n_32_397), .A3(
      multiplier_0_n_32_398));
  DFFR_X1_LVT \multiplier_0_op1_reg[8] (.Q(multiplier_0_op1[8]), .QN(), .CK(
      multiplier_0_n_41), .D(multiplier_0_per_din_msk[8]), .RN(multiplier_0_n_38));
  NAND2_X1_LVT multiplier_0_i_32_76 (.ZN(multiplier_0_n_32_76), .A1(
      multiplier_0_op2_xp[4]), .A2(multiplier_0_op1[8]));
  NAND2_X1_LVT multiplier_0_i_32_92 (.ZN(multiplier_0_n_32_92), .A1(
      multiplier_0_op2_xp[5]), .A2(multiplier_0_op1[7]));
  NOR2_X1_LVT multiplier_0_i_32_366 (.ZN(multiplier_0_n_32_389), .A1(
      multiplier_0_n_32_76), .A2(multiplier_0_n_32_92));
  DFFR_X1_LVT \multiplier_0_op1_reg[9] (.Q(multiplier_0_op1[9]), .QN(), .CK(
      multiplier_0_n_41), .D(multiplier_0_per_din_msk[9]), .RN(multiplier_0_n_38));
  NAND2_X1_LVT multiplier_0_i_32_60 (.ZN(multiplier_0_n_32_60), .A1(
      multiplier_0_op2_xp[3]), .A2(multiplier_0_op1[9]));
  NOR2_X1_LVT multiplier_0_i_32_367 (.ZN(multiplier_0_n_32_390), .A1(
      multiplier_0_n_32_60), .A2(multiplier_0_n_32_92));
  NOR2_X1_LVT multiplier_0_i_32_368 (.ZN(multiplier_0_n_32_391), .A1(
      multiplier_0_n_32_60), .A2(multiplier_0_n_32_76));
  OR3_X1_LVT multiplier_0_i_32_365 (.ZN(multiplier_0_n_32_388), .A1(
      multiplier_0_n_32_389), .A2(multiplier_0_n_32_390), .A3(
      multiplier_0_n_32_391));
  NAND2_X1_LVT multiplier_0_i_32_140 (.ZN(multiplier_0_n_32_140), .A1(
      multiplier_0_op2_xp[8]), .A2(multiplier_0_op1[4]));
  NAND2_X1_LVT multiplier_0_i_32_124 (.ZN(multiplier_0_n_32_124), .A1(
      multiplier_0_op2_xp[7]), .A2(multiplier_0_op1[5]));
  INV_X1_LVT multiplier_0_i_32_358 (.ZN(multiplier_0_n_32_381), .A(
      multiplier_0_n_32_124));
  NAND2_X1_LVT multiplier_0_i_32_357 (.ZN(multiplier_0_n_32_380), .A1(
      multiplier_0_n_32_140), .A2(multiplier_0_n_32_381));
  NAND2_X1_LVT multiplier_0_i_32_108 (.ZN(multiplier_0_n_32_108), .A1(
      multiplier_0_op2_xp[6]), .A2(multiplier_0_op1[6]));
  INV_X1_LVT multiplier_0_i_32_360 (.ZN(multiplier_0_n_32_383), .A(
      multiplier_0_n_32_108));
  NAND2_X1_LVT multiplier_0_i_32_359 (.ZN(multiplier_0_n_32_382), .A1(
      multiplier_0_n_32_140), .A2(multiplier_0_n_32_383));
  OR2_X1_LVT multiplier_0_i_32_361 (.ZN(multiplier_0_n_32_384), .A1(
      multiplier_0_n_32_108), .A2(multiplier_0_n_32_124));
  NAND3_X1_LVT multiplier_0_i_32_356 (.ZN(multiplier_0_n_32_379), .A1(
      multiplier_0_n_32_380), .A2(multiplier_0_n_32_382), .A3(
      multiplier_0_n_32_384));
  FA_X1_LVT multiplier_0_i_32_402 (.CO(multiplier_0_n_32_430), .S(
      multiplier_0_n_32_429), .A(multiplier_0_n_32_395), .B(
      multiplier_0_n_32_388), .CI(multiplier_0_n_32_379));
  NAND2_X1_LVT multiplier_0_i_32_26 (.ZN(multiplier_0_n_32_26), .A1(
      multiplier_0_op2_xp[1]), .A2(multiplier_0_op1[9]));
  NAND2_X1_LVT multiplier_0_i_32_42 (.ZN(multiplier_0_n_32_42), .A1(
      multiplier_0_op2_xp[2]), .A2(multiplier_0_op1[8]));
  NOR2_X1_LVT multiplier_0_i_32_321 (.ZN(multiplier_0_n_32_336), .A1(
      multiplier_0_n_32_26), .A2(multiplier_0_n_32_42));
  NAND2_X1_LVT multiplier_0_i_32_10 (.ZN(multiplier_0_n_32_10), .A1(
      multiplier_0_op2_xp[0]), .A2(multiplier_0_op1[10]));
  NOR2_X1_LVT multiplier_0_i_32_322 (.ZN(multiplier_0_n_32_337), .A1(
      multiplier_0_n_32_10), .A2(multiplier_0_n_32_42));
  NOR2_X1_LVT multiplier_0_i_32_323 (.ZN(multiplier_0_n_32_338), .A1(
      multiplier_0_n_32_10), .A2(multiplier_0_n_32_26));
  OR3_X1_LVT multiplier_0_i_32_320 (.ZN(multiplier_0_n_32_335), .A1(
      multiplier_0_n_32_336), .A2(multiplier_0_n_32_337), .A3(
      multiplier_0_n_32_338));
  NAND2_X1_LVT multiplier_0_i_32_74 (.ZN(multiplier_0_n_32_74), .A1(
      multiplier_0_op2_xp[4]), .A2(multiplier_0_op1[6]));
  NAND2_X1_LVT multiplier_0_i_32_90 (.ZN(multiplier_0_n_32_90), .A1(
      multiplier_0_op2_xp[5]), .A2(multiplier_0_op1[5]));
  NOR2_X1_LVT multiplier_0_i_32_314 (.ZN(multiplier_0_n_32_329), .A1(
      multiplier_0_n_32_74), .A2(multiplier_0_n_32_90));
  NAND2_X1_LVT multiplier_0_i_32_58 (.ZN(multiplier_0_n_32_58), .A1(
      multiplier_0_op2_xp[3]), .A2(multiplier_0_op1[7]));
  NOR2_X1_LVT multiplier_0_i_32_315 (.ZN(multiplier_0_n_32_330), .A1(
      multiplier_0_n_32_58), .A2(multiplier_0_n_32_90));
  NOR2_X1_LVT multiplier_0_i_32_316 (.ZN(multiplier_0_n_32_331), .A1(
      multiplier_0_n_32_58), .A2(multiplier_0_n_32_74));
  OR3_X1_LVT multiplier_0_i_32_313 (.ZN(multiplier_0_n_32_328), .A1(
      multiplier_0_n_32_329), .A2(multiplier_0_n_32_330), .A3(
      multiplier_0_n_32_331));
  NAND2_X1_LVT multiplier_0_i_32_138 (.ZN(multiplier_0_n_32_138), .A1(
      multiplier_0_op2_xp[8]), .A2(multiplier_0_op1[2]));
  NAND2_X1_LVT multiplier_0_i_32_122 (.ZN(multiplier_0_n_32_122), .A1(
      multiplier_0_op2_xp[7]), .A2(multiplier_0_op1[3]));
  INV_X1_LVT multiplier_0_i_32_306 (.ZN(multiplier_0_n_32_321), .A(
      multiplier_0_n_32_122));
  NAND2_X1_LVT multiplier_0_i_32_305 (.ZN(multiplier_0_n_32_320), .A1(
      multiplier_0_n_32_138), .A2(multiplier_0_n_32_321));
  NAND2_X1_LVT multiplier_0_i_32_106 (.ZN(multiplier_0_n_32_106), .A1(
      multiplier_0_op2_xp[6]), .A2(multiplier_0_op1[4]));
  INV_X1_LVT multiplier_0_i_32_308 (.ZN(multiplier_0_n_32_323), .A(
      multiplier_0_n_32_106));
  NAND2_X1_LVT multiplier_0_i_32_307 (.ZN(multiplier_0_n_32_322), .A1(
      multiplier_0_n_32_138), .A2(multiplier_0_n_32_323));
  OR2_X1_LVT multiplier_0_i_32_309 (.ZN(multiplier_0_n_32_324), .A1(
      multiplier_0_n_32_106), .A2(multiplier_0_n_32_122));
  NAND3_X1_LVT multiplier_0_i_32_304 (.ZN(multiplier_0_n_32_319), .A1(
      multiplier_0_n_32_320), .A2(multiplier_0_n_32_322), .A3(
      multiplier_0_n_32_324));
  FA_X1_LVT multiplier_0_i_32_350 (.CO(multiplier_0_n_32_370), .S(
      multiplier_0_n_32_369), .A(multiplier_0_n_32_335), .B(
      multiplier_0_n_32_328), .CI(multiplier_0_n_32_319));
  XNOR2_X1_LVT multiplier_0_i_32_369 (.ZN(multiplier_0_n_32_392), .A(
      multiplier_0_n_32_44), .B(multiplier_0_n_32_28));
  XNOR2_X1_LVT multiplier_0_i_32_370 (.ZN(multiplier_0_n_32_393), .A(
      multiplier_0_n_32_392), .B(multiplier_0_n_32_12));
  INV_X1_LVT multiplier_0_i_32_371 (.ZN(multiplier_0_n_32_394), .A(
      multiplier_0_n_32_393));
  XNOR2_X1_LVT multiplier_0_i_32_362 (.ZN(multiplier_0_n_32_385), .A(
      multiplier_0_n_32_92), .B(multiplier_0_n_32_76));
  XNOR2_X1_LVT multiplier_0_i_32_363 (.ZN(multiplier_0_n_32_386), .A(
      multiplier_0_n_32_385), .B(multiplier_0_n_32_60));
  INV_X1_LVT multiplier_0_i_32_364 (.ZN(multiplier_0_n_32_387), .A(
      multiplier_0_n_32_386));
  FA_X1_LVT multiplier_0_i_32_377 (.CO(multiplier_0_n_32_402), .S(
      multiplier_0_n_32_401), .A(multiplier_0_n_32_370), .B(
      multiplier_0_n_32_394), .CI(multiplier_0_n_32_387));
  FA_X1_LVT multiplier_0_i_32_404 (.CO(multiplier_0_n_32_434), .S(
      multiplier_0_n_32_433), .A(multiplier_0_n_32_408), .B(
      multiplier_0_n_32_429), .CI(multiplier_0_n_32_402));
  NAND2_X1_LVT multiplier_0_i_32_46 (.ZN(multiplier_0_n_32_46), .A1(
      multiplier_0_op2_xp[2]), .A2(multiplier_0_op1[12]));
  DFFR_X1_LVT \multiplier_0_op1_reg[13] (.Q(multiplier_0_op1[13]), .QN(), .CK(
      multiplier_0_n_41), .D(multiplier_0_per_din_msk[13]), .RN(
      multiplier_0_n_38));
  NAND2_X1_LVT multiplier_0_i_32_30 (.ZN(multiplier_0_n_32_30), .A1(
      multiplier_0_op2_xp[1]), .A2(multiplier_0_op1[13]));
  XNOR2_X1_LVT multiplier_0_i_32_421 (.ZN(multiplier_0_n_32_452), .A(
      multiplier_0_n_32_46), .B(multiplier_0_n_32_30));
  DFFR_X1_LVT \multiplier_0_op1_reg[14] (.Q(multiplier_0_op1[14]), .QN(), .CK(
      multiplier_0_n_41), .D(multiplier_0_per_din_msk[14]), .RN(
      multiplier_0_n_38));
  NAND2_X1_LVT multiplier_0_i_32_14 (.ZN(multiplier_0_n_32_14), .A1(
      multiplier_0_op2_xp[0]), .A2(multiplier_0_op1[14]));
  XNOR2_X1_LVT multiplier_0_i_32_422 (.ZN(multiplier_0_n_32_453), .A(
      multiplier_0_n_32_452), .B(multiplier_0_n_32_14));
  INV_X1_LVT multiplier_0_i_32_423 (.ZN(multiplier_0_n_32_454), .A(
      multiplier_0_n_32_453));
  NAND2_X1_LVT multiplier_0_i_32_94 (.ZN(multiplier_0_n_32_94), .A1(
      multiplier_0_op2_xp[5]), .A2(multiplier_0_op1[9]));
  NAND2_X1_LVT multiplier_0_i_32_78 (.ZN(multiplier_0_n_32_78), .A1(
      multiplier_0_op2_xp[4]), .A2(multiplier_0_op1[10]));
  XNOR2_X1_LVT multiplier_0_i_32_414 (.ZN(multiplier_0_n_32_445), .A(
      multiplier_0_n_32_94), .B(multiplier_0_n_32_78));
  NAND2_X1_LVT multiplier_0_i_32_62 (.ZN(multiplier_0_n_32_62), .A1(
      multiplier_0_op2_xp[3]), .A2(multiplier_0_op1[11]));
  XNOR2_X1_LVT multiplier_0_i_32_415 (.ZN(multiplier_0_n_32_446), .A(
      multiplier_0_n_32_445), .B(multiplier_0_n_32_62));
  INV_X1_LVT multiplier_0_i_32_416 (.ZN(multiplier_0_n_32_447), .A(
      multiplier_0_n_32_446));
  FA_X1_LVT multiplier_0_i_32_429 (.CO(multiplier_0_n_32_462), .S(
      multiplier_0_n_32_461), .A(multiplier_0_n_32_430), .B(
      multiplier_0_n_32_454), .CI(multiplier_0_n_32_447));
  NAND2_X1_LVT multiplier_0_i_32_142 (.ZN(multiplier_0_n_32_142), .A1(
      multiplier_0_op2_xp[8]), .A2(multiplier_0_op1[6]));
  NAND2_X1_LVT multiplier_0_i_32_126 (.ZN(multiplier_0_n_32_126), .A1(
      multiplier_0_op2_xp[7]), .A2(multiplier_0_op1[7]));
  XNOR2_X1_LVT multiplier_0_i_32_406 (.ZN(multiplier_0_n_32_437), .A(
      multiplier_0_n_32_142), .B(multiplier_0_n_32_126));
  NAND2_X1_LVT multiplier_0_i_32_110 (.ZN(multiplier_0_n_32_110), .A1(
      multiplier_0_op2_xp[6]), .A2(multiplier_0_op1[8]));
  XNOR2_X1_LVT multiplier_0_i_32_407 (.ZN(multiplier_0_n_32_438), .A(
      multiplier_0_n_32_437), .B(multiplier_0_n_32_110));
  NAND2_X1_LVT multiplier_0_i_32_29 (.ZN(multiplier_0_n_32_29), .A1(
      multiplier_0_op2_xp[1]), .A2(multiplier_0_op1[12]));
  NAND2_X1_LVT multiplier_0_i_32_45 (.ZN(multiplier_0_n_32_45), .A1(
      multiplier_0_op2_xp[2]), .A2(multiplier_0_op1[11]));
  NOR2_X1_LVT multiplier_0_i_32_399 (.ZN(multiplier_0_n_32_426), .A1(
      multiplier_0_n_32_29), .A2(multiplier_0_n_32_45));
  NAND2_X1_LVT multiplier_0_i_32_13 (.ZN(multiplier_0_n_32_13), .A1(
      multiplier_0_op2_xp[0]), .A2(multiplier_0_op1[13]));
  NOR2_X1_LVT multiplier_0_i_32_400 (.ZN(multiplier_0_n_32_427), .A1(
      multiplier_0_n_32_13), .A2(multiplier_0_n_32_45));
  NOR2_X1_LVT multiplier_0_i_32_401 (.ZN(multiplier_0_n_32_428), .A1(
      multiplier_0_n_32_13), .A2(multiplier_0_n_32_29));
  OR3_X1_LVT multiplier_0_i_32_398 (.ZN(multiplier_0_n_32_425), .A1(
      multiplier_0_n_32_426), .A2(multiplier_0_n_32_427), .A3(
      multiplier_0_n_32_428));
  NAND2_X1_LVT multiplier_0_i_32_77 (.ZN(multiplier_0_n_32_77), .A1(
      multiplier_0_op2_xp[4]), .A2(multiplier_0_op1[9]));
  NAND2_X1_LVT multiplier_0_i_32_93 (.ZN(multiplier_0_n_32_93), .A1(
      multiplier_0_op2_xp[5]), .A2(multiplier_0_op1[8]));
  NOR2_X1_LVT multiplier_0_i_32_392 (.ZN(multiplier_0_n_32_419), .A1(
      multiplier_0_n_32_77), .A2(multiplier_0_n_32_93));
  NAND2_X1_LVT multiplier_0_i_32_61 (.ZN(multiplier_0_n_32_61), .A1(
      multiplier_0_op2_xp[3]), .A2(multiplier_0_op1[10]));
  NOR2_X1_LVT multiplier_0_i_32_393 (.ZN(multiplier_0_n_32_420), .A1(
      multiplier_0_n_32_61), .A2(multiplier_0_n_32_93));
  NOR2_X1_LVT multiplier_0_i_32_394 (.ZN(multiplier_0_n_32_421), .A1(
      multiplier_0_n_32_61), .A2(multiplier_0_n_32_77));
  OR3_X1_LVT multiplier_0_i_32_391 (.ZN(multiplier_0_n_32_418), .A1(
      multiplier_0_n_32_419), .A2(multiplier_0_n_32_420), .A3(
      multiplier_0_n_32_421));
  INV_X1_LVT multiplier_0_i_32_384 (.ZN(multiplier_0_n_32_411), .A(
      multiplier_0_n_32_125));
  NAND2_X1_LVT multiplier_0_i_32_383 (.ZN(multiplier_0_n_32_410), .A1(
      multiplier_0_n_32_141), .A2(multiplier_0_n_32_411));
  INV_X1_LVT multiplier_0_i_32_386 (.ZN(multiplier_0_n_32_413), .A(
      multiplier_0_n_32_109));
  NAND2_X1_LVT multiplier_0_i_32_385 (.ZN(multiplier_0_n_32_412), .A1(
      multiplier_0_n_32_141), .A2(multiplier_0_n_32_413));
  OR2_X1_LVT multiplier_0_i_32_387 (.ZN(multiplier_0_n_32_414), .A1(
      multiplier_0_n_32_109), .A2(multiplier_0_n_32_125));
  NAND3_X1_LVT multiplier_0_i_32_382 (.ZN(multiplier_0_n_32_409), .A1(
      multiplier_0_n_32_410), .A2(multiplier_0_n_32_412), .A3(
      multiplier_0_n_32_414));
  FA_X1_LVT multiplier_0_i_32_428 (.CO(multiplier_0_n_32_460), .S(
      multiplier_0_n_32_459), .A(multiplier_0_n_32_425), .B(
      multiplier_0_n_32_418), .CI(multiplier_0_n_32_409));
  NAND2_X1_LVT multiplier_0_i_32_27 (.ZN(multiplier_0_n_32_27), .A1(
      multiplier_0_op2_xp[1]), .A2(multiplier_0_op1[10]));
  NAND2_X1_LVT multiplier_0_i_32_43 (.ZN(multiplier_0_n_32_43), .A1(
      multiplier_0_op2_xp[2]), .A2(multiplier_0_op1[9]));
  NOR2_X1_LVT multiplier_0_i_32_347 (.ZN(multiplier_0_n_32_366), .A1(
      multiplier_0_n_32_27), .A2(multiplier_0_n_32_43));
  NAND2_X1_LVT multiplier_0_i_32_11 (.ZN(multiplier_0_n_32_11), .A1(
      multiplier_0_op2_xp[0]), .A2(multiplier_0_op1[11]));
  NOR2_X1_LVT multiplier_0_i_32_348 (.ZN(multiplier_0_n_32_367), .A1(
      multiplier_0_n_32_11), .A2(multiplier_0_n_32_43));
  NOR2_X1_LVT multiplier_0_i_32_349 (.ZN(multiplier_0_n_32_368), .A1(
      multiplier_0_n_32_11), .A2(multiplier_0_n_32_27));
  OR3_X1_LVT multiplier_0_i_32_346 (.ZN(multiplier_0_n_32_365), .A1(
      multiplier_0_n_32_366), .A2(multiplier_0_n_32_367), .A3(
      multiplier_0_n_32_368));
  NAND2_X1_LVT multiplier_0_i_32_75 (.ZN(multiplier_0_n_32_75), .A1(
      multiplier_0_op2_xp[4]), .A2(multiplier_0_op1[7]));
  NAND2_X1_LVT multiplier_0_i_32_91 (.ZN(multiplier_0_n_32_91), .A1(
      multiplier_0_op2_xp[5]), .A2(multiplier_0_op1[6]));
  NOR2_X1_LVT multiplier_0_i_32_340 (.ZN(multiplier_0_n_32_359), .A1(
      multiplier_0_n_32_75), .A2(multiplier_0_n_32_91));
  NAND2_X1_LVT multiplier_0_i_32_59 (.ZN(multiplier_0_n_32_59), .A1(
      multiplier_0_op2_xp[3]), .A2(multiplier_0_op1[8]));
  NOR2_X1_LVT multiplier_0_i_32_341 (.ZN(multiplier_0_n_32_360), .A1(
      multiplier_0_n_32_59), .A2(multiplier_0_n_32_91));
  NOR2_X1_LVT multiplier_0_i_32_342 (.ZN(multiplier_0_n_32_361), .A1(
      multiplier_0_n_32_59), .A2(multiplier_0_n_32_75));
  OR3_X1_LVT multiplier_0_i_32_339 (.ZN(multiplier_0_n_32_358), .A1(
      multiplier_0_n_32_359), .A2(multiplier_0_n_32_360), .A3(
      multiplier_0_n_32_361));
  NAND2_X1_LVT multiplier_0_i_32_139 (.ZN(multiplier_0_n_32_139), .A1(
      multiplier_0_op2_xp[8]), .A2(multiplier_0_op1[3]));
  NAND2_X1_LVT multiplier_0_i_32_123 (.ZN(multiplier_0_n_32_123), .A1(
      multiplier_0_op2_xp[7]), .A2(multiplier_0_op1[4]));
  INV_X1_LVT multiplier_0_i_32_332 (.ZN(multiplier_0_n_32_351), .A(
      multiplier_0_n_32_123));
  NAND2_X1_LVT multiplier_0_i_32_331 (.ZN(multiplier_0_n_32_350), .A1(
      multiplier_0_n_32_139), .A2(multiplier_0_n_32_351));
  NAND2_X1_LVT multiplier_0_i_32_107 (.ZN(multiplier_0_n_32_107), .A1(
      multiplier_0_op2_xp[6]), .A2(multiplier_0_op1[5]));
  INV_X1_LVT multiplier_0_i_32_334 (.ZN(multiplier_0_n_32_353), .A(
      multiplier_0_n_32_107));
  NAND2_X1_LVT multiplier_0_i_32_333 (.ZN(multiplier_0_n_32_352), .A1(
      multiplier_0_n_32_139), .A2(multiplier_0_n_32_353));
  OR2_X1_LVT multiplier_0_i_32_335 (.ZN(multiplier_0_n_32_354), .A1(
      multiplier_0_n_32_107), .A2(multiplier_0_n_32_123));
  NAND3_X1_LVT multiplier_0_i_32_330 (.ZN(multiplier_0_n_32_349), .A1(
      multiplier_0_n_32_350), .A2(multiplier_0_n_32_352), .A3(
      multiplier_0_n_32_354));
  FA_X1_LVT multiplier_0_i_32_376 (.CO(multiplier_0_n_32_400), .S(
      multiplier_0_n_32_399), .A(multiplier_0_n_32_365), .B(
      multiplier_0_n_32_358), .CI(multiplier_0_n_32_349));
  XNOR2_X1_LVT multiplier_0_i_32_395 (.ZN(multiplier_0_n_32_422), .A(
      multiplier_0_n_32_45), .B(multiplier_0_n_32_29));
  XNOR2_X1_LVT multiplier_0_i_32_396 (.ZN(multiplier_0_n_32_423), .A(
      multiplier_0_n_32_422), .B(multiplier_0_n_32_13));
  INV_X1_LVT multiplier_0_i_32_397 (.ZN(multiplier_0_n_32_424), .A(
      multiplier_0_n_32_423));
  XNOR2_X1_LVT multiplier_0_i_32_388 (.ZN(multiplier_0_n_32_415), .A(
      multiplier_0_n_32_93), .B(multiplier_0_n_32_77));
  XNOR2_X1_LVT multiplier_0_i_32_389 (.ZN(multiplier_0_n_32_416), .A(
      multiplier_0_n_32_415), .B(multiplier_0_n_32_61));
  INV_X1_LVT multiplier_0_i_32_390 (.ZN(multiplier_0_n_32_417), .A(
      multiplier_0_n_32_416));
  FA_X1_LVT multiplier_0_i_32_403 (.CO(multiplier_0_n_32_432), .S(
      multiplier_0_n_32_431), .A(multiplier_0_n_32_400), .B(
      multiplier_0_n_32_424), .CI(multiplier_0_n_32_417));
  FA_X1_LVT multiplier_0_i_32_430 (.CO(multiplier_0_n_32_464), .S(
      multiplier_0_n_32_463), .A(multiplier_0_n_32_438), .B(
      multiplier_0_n_32_459), .CI(multiplier_0_n_32_432));
  FA_X1_LVT multiplier_0_i_32_431 (.CO(multiplier_0_n_32_466), .S(
      multiplier_0_n_32_465), .A(multiplier_0_n_32_434), .B(
      multiplier_0_n_32_461), .CI(multiplier_0_n_32_463));
  NAND2_X1_LVT multiplier_0_i_32_47 (.ZN(multiplier_0_n_32_47), .A1(
      multiplier_0_op2_xp[2]), .A2(multiplier_0_op1[13]));
  NAND2_X1_LVT multiplier_0_i_32_31 (.ZN(multiplier_0_n_32_31), .A1(
      multiplier_0_op2_xp[1]), .A2(multiplier_0_op1[14]));
  XNOR2_X1_LVT multiplier_0_i_32_447 (.ZN(multiplier_0_n_32_482), .A(
      multiplier_0_n_32_47), .B(multiplier_0_n_32_31));
  DFFR_X1_LVT \multiplier_0_op1_reg[15] (.Q(multiplier_0_op1[15]), .QN(), .CK(
      multiplier_0_n_41), .D(multiplier_0_per_din_msk[15]), .RN(
      multiplier_0_n_38));
  NAND2_X1_LVT multiplier_0_i_32_15 (.ZN(multiplier_0_n_32_15), .A1(
      multiplier_0_op2_xp[0]), .A2(multiplier_0_op1[15]));
  XNOR2_X1_LVT multiplier_0_i_32_448 (.ZN(multiplier_0_n_32_483), .A(
      multiplier_0_n_32_482), .B(multiplier_0_n_32_15));
  INV_X1_LVT multiplier_0_i_32_449 (.ZN(multiplier_0_n_32_484), .A(
      multiplier_0_n_32_483));
  NAND2_X1_LVT multiplier_0_i_32_95 (.ZN(multiplier_0_n_32_95), .A1(
      multiplier_0_op2_xp[5]), .A2(multiplier_0_op1[10]));
  NAND2_X1_LVT multiplier_0_i_32_79 (.ZN(multiplier_0_n_32_79), .A1(
      multiplier_0_op2_xp[4]), .A2(multiplier_0_op1[11]));
  XNOR2_X1_LVT multiplier_0_i_32_440 (.ZN(multiplier_0_n_32_475), .A(
      multiplier_0_n_32_95), .B(multiplier_0_n_32_79));
  NAND2_X1_LVT multiplier_0_i_32_63 (.ZN(multiplier_0_n_32_63), .A1(
      multiplier_0_op2_xp[3]), .A2(multiplier_0_op1[12]));
  XNOR2_X1_LVT multiplier_0_i_32_441 (.ZN(multiplier_0_n_32_476), .A(
      multiplier_0_n_32_475), .B(multiplier_0_n_32_63));
  INV_X1_LVT multiplier_0_i_32_442 (.ZN(multiplier_0_n_32_477), .A(
      multiplier_0_n_32_476));
  FA_X1_LVT multiplier_0_i_32_455 (.CO(multiplier_0_n_32_492), .S(
      multiplier_0_n_32_491), .A(multiplier_0_n_32_460), .B(
      multiplier_0_n_32_484), .CI(multiplier_0_n_32_477));
  NAND2_X1_LVT multiplier_0_i_32_143 (.ZN(multiplier_0_n_32_143), .A1(
      multiplier_0_op2_xp[8]), .A2(multiplier_0_op1[7]));
  NAND2_X1_LVT multiplier_0_i_32_127 (.ZN(multiplier_0_n_32_127), .A1(
      multiplier_0_op2_xp[7]), .A2(multiplier_0_op1[8]));
  XNOR2_X1_LVT multiplier_0_i_32_432 (.ZN(multiplier_0_n_32_467), .A(
      multiplier_0_n_32_143), .B(multiplier_0_n_32_127));
  NAND2_X1_LVT multiplier_0_i_32_111 (.ZN(multiplier_0_n_32_111), .A1(
      multiplier_0_op2_xp[6]), .A2(multiplier_0_op1[9]));
  XNOR2_X1_LVT multiplier_0_i_32_433 (.ZN(multiplier_0_n_32_468), .A(
      multiplier_0_n_32_467), .B(multiplier_0_n_32_111));
  NOR2_X1_LVT multiplier_0_i_32_425 (.ZN(multiplier_0_n_32_456), .A1(
      multiplier_0_n_32_30), .A2(multiplier_0_n_32_46));
  NOR2_X1_LVT multiplier_0_i_32_426 (.ZN(multiplier_0_n_32_457), .A1(
      multiplier_0_n_32_14), .A2(multiplier_0_n_32_46));
  NOR2_X1_LVT multiplier_0_i_32_427 (.ZN(multiplier_0_n_32_458), .A1(
      multiplier_0_n_32_14), .A2(multiplier_0_n_32_30));
  OR3_X1_LVT multiplier_0_i_32_424 (.ZN(multiplier_0_n_32_455), .A1(
      multiplier_0_n_32_456), .A2(multiplier_0_n_32_457), .A3(
      multiplier_0_n_32_458));
  NOR2_X1_LVT multiplier_0_i_32_418 (.ZN(multiplier_0_n_32_449), .A1(
      multiplier_0_n_32_78), .A2(multiplier_0_n_32_94));
  NOR2_X1_LVT multiplier_0_i_32_419 (.ZN(multiplier_0_n_32_450), .A1(
      multiplier_0_n_32_62), .A2(multiplier_0_n_32_94));
  NOR2_X1_LVT multiplier_0_i_32_420 (.ZN(multiplier_0_n_32_451), .A1(
      multiplier_0_n_32_62), .A2(multiplier_0_n_32_78));
  OR3_X1_LVT multiplier_0_i_32_417 (.ZN(multiplier_0_n_32_448), .A1(
      multiplier_0_n_32_449), .A2(multiplier_0_n_32_450), .A3(
      multiplier_0_n_32_451));
  INV_X1_LVT multiplier_0_i_32_410 (.ZN(multiplier_0_n_32_441), .A(
      multiplier_0_n_32_126));
  NAND2_X1_LVT multiplier_0_i_32_409 (.ZN(multiplier_0_n_32_440), .A1(
      multiplier_0_n_32_142), .A2(multiplier_0_n_32_441));
  INV_X1_LVT multiplier_0_i_32_412 (.ZN(multiplier_0_n_32_443), .A(
      multiplier_0_n_32_110));
  NAND2_X1_LVT multiplier_0_i_32_411 (.ZN(multiplier_0_n_32_442), .A1(
      multiplier_0_n_32_142), .A2(multiplier_0_n_32_443));
  OR2_X1_LVT multiplier_0_i_32_413 (.ZN(multiplier_0_n_32_444), .A1(
      multiplier_0_n_32_110), .A2(multiplier_0_n_32_126));
  NAND3_X1_LVT multiplier_0_i_32_408 (.ZN(multiplier_0_n_32_439), .A1(
      multiplier_0_n_32_440), .A2(multiplier_0_n_32_442), .A3(
      multiplier_0_n_32_444));
  FA_X1_LVT multiplier_0_i_32_454 (.CO(multiplier_0_n_32_490), .S(
      multiplier_0_n_32_489), .A(multiplier_0_n_32_455), .B(
      multiplier_0_n_32_448), .CI(multiplier_0_n_32_439));
  FA_X1_LVT multiplier_0_i_32_456 (.CO(multiplier_0_n_32_494), .S(
      multiplier_0_n_32_493), .A(multiplier_0_n_32_468), .B(
      multiplier_0_n_32_489), .CI(multiplier_0_n_32_462));
  FA_X1_LVT multiplier_0_i_32_457 (.CO(multiplier_0_n_32_496), .S(
      multiplier_0_n_32_495), .A(multiplier_0_n_32_464), .B(
      multiplier_0_n_32_491), .CI(multiplier_0_n_32_493));
  XNOR2_X1_LVT multiplier_0_i_32_354 (.ZN(multiplier_0_n_32_377), .A(
      multiplier_0_n_32_140), .B(multiplier_0_n_32_124));
  XNOR2_X1_LVT multiplier_0_i_32_355 (.ZN(multiplier_0_n_32_378), .A(
      multiplier_0_n_32_377), .B(multiplier_0_n_32_108));
  NAND2_X1_LVT multiplier_0_i_32_25 (.ZN(multiplier_0_n_32_25), .A1(
      multiplier_0_op2_xp[1]), .A2(multiplier_0_op1[8]));
  NAND2_X1_LVT multiplier_0_i_32_41 (.ZN(multiplier_0_n_32_41), .A1(
      multiplier_0_op2_xp[2]), .A2(multiplier_0_op1[7]));
  NOR2_X1_LVT multiplier_0_i_32_295 (.ZN(multiplier_0_n_32_306), .A1(
      multiplier_0_n_32_25), .A2(multiplier_0_n_32_41));
  NAND2_X1_LVT multiplier_0_i_32_9 (.ZN(multiplier_0_n_32_9), .A1(
      multiplier_0_op2_xp[0]), .A2(multiplier_0_op1[9]));
  NOR2_X1_LVT multiplier_0_i_32_296 (.ZN(multiplier_0_n_32_307), .A1(
      multiplier_0_n_32_9), .A2(multiplier_0_n_32_41));
  NOR2_X1_LVT multiplier_0_i_32_297 (.ZN(multiplier_0_n_32_308), .A1(
      multiplier_0_n_32_9), .A2(multiplier_0_n_32_25));
  OR3_X1_LVT multiplier_0_i_32_294 (.ZN(multiplier_0_n_32_305), .A1(
      multiplier_0_n_32_306), .A2(multiplier_0_n_32_307), .A3(
      multiplier_0_n_32_308));
  NAND2_X1_LVT multiplier_0_i_32_73 (.ZN(multiplier_0_n_32_73), .A1(
      multiplier_0_op2_xp[4]), .A2(multiplier_0_op1[5]));
  NAND2_X1_LVT multiplier_0_i_32_89 (.ZN(multiplier_0_n_32_89), .A1(
      multiplier_0_op2_xp[5]), .A2(multiplier_0_op1[4]));
  NOR2_X1_LVT multiplier_0_i_32_288 (.ZN(multiplier_0_n_32_299), .A1(
      multiplier_0_n_32_73), .A2(multiplier_0_n_32_89));
  NAND2_X1_LVT multiplier_0_i_32_57 (.ZN(multiplier_0_n_32_57), .A1(
      multiplier_0_op2_xp[3]), .A2(multiplier_0_op1[6]));
  NOR2_X1_LVT multiplier_0_i_32_289 (.ZN(multiplier_0_n_32_300), .A1(
      multiplier_0_n_32_57), .A2(multiplier_0_n_32_89));
  NOR2_X1_LVT multiplier_0_i_32_290 (.ZN(multiplier_0_n_32_301), .A1(
      multiplier_0_n_32_57), .A2(multiplier_0_n_32_73));
  OR3_X1_LVT multiplier_0_i_32_287 (.ZN(multiplier_0_n_32_298), .A1(
      multiplier_0_n_32_299), .A2(multiplier_0_n_32_300), .A3(
      multiplier_0_n_32_301));
  NAND2_X1_LVT multiplier_0_i_32_137 (.ZN(multiplier_0_n_32_137), .A1(
      multiplier_0_op2_xp[8]), .A2(multiplier_0_op1[1]));
  NAND2_X1_LVT multiplier_0_i_32_121 (.ZN(multiplier_0_n_32_121), .A1(
      multiplier_0_op2_xp[7]), .A2(multiplier_0_op1[2]));
  INV_X1_LVT multiplier_0_i_32_280 (.ZN(multiplier_0_n_32_291), .A(
      multiplier_0_n_32_121));
  NAND2_X1_LVT multiplier_0_i_32_279 (.ZN(multiplier_0_n_32_290), .A1(
      multiplier_0_n_32_137), .A2(multiplier_0_n_32_291));
  NAND2_X1_LVT multiplier_0_i_32_105 (.ZN(multiplier_0_n_32_105), .A1(
      multiplier_0_op2_xp[6]), .A2(multiplier_0_op1[3]));
  INV_X1_LVT multiplier_0_i_32_282 (.ZN(multiplier_0_n_32_293), .A(
      multiplier_0_n_32_105));
  NAND2_X1_LVT multiplier_0_i_32_281 (.ZN(multiplier_0_n_32_292), .A1(
      multiplier_0_n_32_137), .A2(multiplier_0_n_32_293));
  OR2_X1_LVT multiplier_0_i_32_283 (.ZN(multiplier_0_n_32_294), .A1(
      multiplier_0_n_32_105), .A2(multiplier_0_n_32_121));
  NAND3_X1_LVT multiplier_0_i_32_278 (.ZN(multiplier_0_n_32_289), .A1(
      multiplier_0_n_32_290), .A2(multiplier_0_n_32_292), .A3(
      multiplier_0_n_32_294));
  FA_X1_LVT multiplier_0_i_32_324 (.CO(multiplier_0_n_32_340), .S(
      multiplier_0_n_32_339), .A(multiplier_0_n_32_305), .B(
      multiplier_0_n_32_298), .CI(multiplier_0_n_32_289));
  XNOR2_X1_LVT multiplier_0_i_32_343 (.ZN(multiplier_0_n_32_362), .A(
      multiplier_0_n_32_43), .B(multiplier_0_n_32_27));
  XNOR2_X1_LVT multiplier_0_i_32_344 (.ZN(multiplier_0_n_32_363), .A(
      multiplier_0_n_32_362), .B(multiplier_0_n_32_11));
  INV_X1_LVT multiplier_0_i_32_345 (.ZN(multiplier_0_n_32_364), .A(
      multiplier_0_n_32_363));
  XNOR2_X1_LVT multiplier_0_i_32_336 (.ZN(multiplier_0_n_32_355), .A(
      multiplier_0_n_32_91), .B(multiplier_0_n_32_75));
  XNOR2_X1_LVT multiplier_0_i_32_337 (.ZN(multiplier_0_n_32_356), .A(
      multiplier_0_n_32_355), .B(multiplier_0_n_32_59));
  INV_X1_LVT multiplier_0_i_32_338 (.ZN(multiplier_0_n_32_357), .A(
      multiplier_0_n_32_356));
  FA_X1_LVT multiplier_0_i_32_351 (.CO(multiplier_0_n_32_372), .S(
      multiplier_0_n_32_371), .A(multiplier_0_n_32_340), .B(
      multiplier_0_n_32_364), .CI(multiplier_0_n_32_357));
  FA_X1_LVT multiplier_0_i_32_378 (.CO(multiplier_0_n_32_404), .S(
      multiplier_0_n_32_403), .A(multiplier_0_n_32_378), .B(
      multiplier_0_n_32_399), .CI(multiplier_0_n_32_372));
  FA_X1_LVT multiplier_0_i_32_405 (.CO(multiplier_0_n_32_436), .S(
      multiplier_0_n_32_435), .A(multiplier_0_n_32_404), .B(
      multiplier_0_n_32_431), .CI(multiplier_0_n_32_433));
  XNOR2_X1_LVT multiplier_0_i_32_328 (.ZN(multiplier_0_n_32_347), .A(
      multiplier_0_n_32_139), .B(multiplier_0_n_32_123));
  XNOR2_X1_LVT multiplier_0_i_32_329 (.ZN(multiplier_0_n_32_348), .A(
      multiplier_0_n_32_347), .B(multiplier_0_n_32_107));
  NAND2_X1_LVT multiplier_0_i_32_40 (.ZN(multiplier_0_n_32_40), .A1(
      multiplier_0_op2_xp[2]), .A2(multiplier_0_op1[6]));
  NAND2_X1_LVT multiplier_0_i_32_56 (.ZN(multiplier_0_n_32_56), .A1(
      multiplier_0_op2_xp[3]), .A2(multiplier_0_op1[5]));
  NOR2_X1_LVT multiplier_0_i_32_262 (.ZN(multiplier_0_n_32_270), .A1(
      multiplier_0_n_32_40), .A2(multiplier_0_n_32_56));
  NAND2_X1_LVT multiplier_0_i_32_24 (.ZN(multiplier_0_n_32_24), .A1(
      multiplier_0_op2_xp[1]), .A2(multiplier_0_op1[7]));
  NOR2_X1_LVT multiplier_0_i_32_263 (.ZN(multiplier_0_n_32_271), .A1(
      multiplier_0_n_32_24), .A2(multiplier_0_n_32_56));
  NOR2_X1_LVT multiplier_0_i_32_264 (.ZN(multiplier_0_n_32_272), .A1(
      multiplier_0_n_32_24), .A2(multiplier_0_n_32_40));
  OR3_X1_LVT multiplier_0_i_32_261 (.ZN(multiplier_0_n_32_269), .A1(
      multiplier_0_n_32_270), .A2(multiplier_0_n_32_271), .A3(
      multiplier_0_n_32_272));
  NAND2_X1_LVT multiplier_0_i_32_88 (.ZN(multiplier_0_n_32_88), .A1(
      multiplier_0_op2_xp[5]), .A2(multiplier_0_op1[3]));
  NAND2_X1_LVT multiplier_0_i_32_104 (.ZN(multiplier_0_n_32_104), .A1(
      multiplier_0_op2_xp[6]), .A2(multiplier_0_op1[2]));
  NOR2_X1_LVT multiplier_0_i_32_255 (.ZN(multiplier_0_n_32_263), .A1(
      multiplier_0_n_32_88), .A2(multiplier_0_n_32_104));
  NAND2_X1_LVT multiplier_0_i_32_72 (.ZN(multiplier_0_n_32_72), .A1(
      multiplier_0_op2_xp[4]), .A2(multiplier_0_op1[4]));
  NOR2_X1_LVT multiplier_0_i_32_256 (.ZN(multiplier_0_n_32_264), .A1(
      multiplier_0_n_32_72), .A2(multiplier_0_n_32_104));
  NOR2_X1_LVT multiplier_0_i_32_257 (.ZN(multiplier_0_n_32_265), .A1(
      multiplier_0_n_32_72), .A2(multiplier_0_n_32_88));
  OR3_X1_LVT multiplier_0_i_32_254 (.ZN(multiplier_0_n_32_262), .A1(
      multiplier_0_n_32_263), .A2(multiplier_0_n_32_264), .A3(
      multiplier_0_n_32_265));
  NAND2_X1_LVT multiplier_0_i_32_120 (.ZN(multiplier_0_n_32_120), .A1(
      multiplier_0_op2_xp[7]), .A2(multiplier_0_op1[1]));
  NAND2_X1_LVT multiplier_0_i_32_136 (.ZN(multiplier_0_n_32_136), .A1(
      multiplier_0_op2_xp[8]), .A2(multiplier_0_op1[0]));
  INV_X1_LVT multiplier_0_i_32_250 (.ZN(multiplier_0_n_32_258), .A(
      multiplier_0_n_32_136));
  NAND2_X1_LVT multiplier_0_i_32_249 (.ZN(multiplier_0_n_32_257), .A1(
      multiplier_0_n_32_120), .A2(multiplier_0_n_32_258));
  FA_X1_LVT multiplier_0_i_32_298 (.CO(multiplier_0_n_32_310), .S(
      multiplier_0_n_32_309), .A(multiplier_0_n_32_269), .B(
      multiplier_0_n_32_262), .CI(multiplier_0_n_32_257));
  XNOR2_X1_LVT multiplier_0_i_32_317 (.ZN(multiplier_0_n_32_332), .A(
      multiplier_0_n_32_42), .B(multiplier_0_n_32_26));
  XNOR2_X1_LVT multiplier_0_i_32_318 (.ZN(multiplier_0_n_32_333), .A(
      multiplier_0_n_32_332), .B(multiplier_0_n_32_10));
  INV_X1_LVT multiplier_0_i_32_319 (.ZN(multiplier_0_n_32_334), .A(
      multiplier_0_n_32_333));
  XNOR2_X1_LVT multiplier_0_i_32_310 (.ZN(multiplier_0_n_32_325), .A(
      multiplier_0_n_32_90), .B(multiplier_0_n_32_74));
  XNOR2_X1_LVT multiplier_0_i_32_311 (.ZN(multiplier_0_n_32_326), .A(
      multiplier_0_n_32_325), .B(multiplier_0_n_32_58));
  INV_X1_LVT multiplier_0_i_32_312 (.ZN(multiplier_0_n_32_327), .A(
      multiplier_0_n_32_326));
  FA_X1_LVT multiplier_0_i_32_325 (.CO(multiplier_0_n_32_342), .S(
      multiplier_0_n_32_341), .A(multiplier_0_n_32_310), .B(
      multiplier_0_n_32_334), .CI(multiplier_0_n_32_327));
  FA_X1_LVT multiplier_0_i_32_352 (.CO(multiplier_0_n_32_374), .S(
      multiplier_0_n_32_373), .A(multiplier_0_n_32_348), .B(
      multiplier_0_n_32_369), .CI(multiplier_0_n_32_342));
  FA_X1_LVT multiplier_0_i_32_379 (.CO(multiplier_0_n_32_406), .S(
      multiplier_0_n_32_405), .A(multiplier_0_n_32_374), .B(
      multiplier_0_n_32_401), .CI(multiplier_0_n_32_403));
  XNOR2_X1_LVT multiplier_0_i_32_302 (.ZN(multiplier_0_n_32_317), .A(
      multiplier_0_n_32_138), .B(multiplier_0_n_32_122));
  XNOR2_X1_LVT multiplier_0_i_32_303 (.ZN(multiplier_0_n_32_318), .A(
      multiplier_0_n_32_317), .B(multiplier_0_n_32_106));
  NOR2_X1_LVT multiplier_0_i_32_233 (.ZN(multiplier_0_n_32_238), .A1(
      multiplier_0_n_32_55), .A2(multiplier_0_n_32_71));
  NOR2_X1_LVT multiplier_0_i_32_234 (.ZN(multiplier_0_n_32_239), .A1(
      multiplier_0_n_32_39), .A2(multiplier_0_n_32_71));
  NOR2_X1_LVT multiplier_0_i_32_235 (.ZN(multiplier_0_n_32_240), .A1(
      multiplier_0_n_32_39), .A2(multiplier_0_n_32_55));
  OR3_X1_LVT multiplier_0_i_32_232 (.ZN(multiplier_0_n_32_237), .A1(
      multiplier_0_n_32_238), .A2(multiplier_0_n_32_239), .A3(
      multiplier_0_n_32_240));
  NAND2_X1_LVT multiplier_0_i_32_8 (.ZN(multiplier_0_n_32_8), .A1(
      multiplier_0_op2_xp[0]), .A2(multiplier_0_op1[8]));
  INV_X1_LVT multiplier_0_i_32_270 (.ZN(multiplier_0_n_32_278), .A(
      multiplier_0_n_32_8));
  NAND2_X1_LVT multiplier_0_i_32_269 (.ZN(multiplier_0_n_32_277), .A1(
      multiplier_0_n_32_237), .A2(multiplier_0_n_32_278));
  NOR2_X1_LVT multiplier_0_i_32_226 (.ZN(multiplier_0_n_32_231), .A1(
      multiplier_0_n_32_103), .A2(multiplier_0_n_32_119));
  NOR2_X1_LVT multiplier_0_i_32_227 (.ZN(multiplier_0_n_32_232), .A1(
      multiplier_0_n_32_87), .A2(multiplier_0_n_32_119));
  NOR2_X1_LVT multiplier_0_i_32_228 (.ZN(multiplier_0_n_32_233), .A1(
      multiplier_0_n_32_87), .A2(multiplier_0_n_32_103));
  OR3_X1_LVT multiplier_0_i_32_225 (.ZN(multiplier_0_n_32_230), .A1(
      multiplier_0_n_32_231), .A2(multiplier_0_n_32_232), .A3(
      multiplier_0_n_32_233));
  NAND2_X1_LVT multiplier_0_i_32_271 (.ZN(multiplier_0_n_32_279), .A1(
      multiplier_0_n_32_230), .A2(multiplier_0_n_32_278));
  NAND2_X1_LVT multiplier_0_i_32_272 (.ZN(multiplier_0_n_32_280), .A1(
      multiplier_0_n_32_230), .A2(multiplier_0_n_32_237));
  NAND3_X1_LVT multiplier_0_i_32_268 (.ZN(multiplier_0_n_32_276), .A1(
      multiplier_0_n_32_277), .A2(multiplier_0_n_32_279), .A3(
      multiplier_0_n_32_280));
  XNOR2_X1_LVT multiplier_0_i_32_291 (.ZN(multiplier_0_n_32_302), .A(
      multiplier_0_n_32_41), .B(multiplier_0_n_32_25));
  XNOR2_X1_LVT multiplier_0_i_32_292 (.ZN(multiplier_0_n_32_303), .A(
      multiplier_0_n_32_302), .B(multiplier_0_n_32_9));
  INV_X1_LVT multiplier_0_i_32_293 (.ZN(multiplier_0_n_32_304), .A(
      multiplier_0_n_32_303));
  XNOR2_X1_LVT multiplier_0_i_32_284 (.ZN(multiplier_0_n_32_295), .A(
      multiplier_0_n_32_89), .B(multiplier_0_n_32_73));
  XNOR2_X1_LVT multiplier_0_i_32_285 (.ZN(multiplier_0_n_32_296), .A(
      multiplier_0_n_32_295), .B(multiplier_0_n_32_57));
  INV_X1_LVT multiplier_0_i_32_286 (.ZN(multiplier_0_n_32_297), .A(
      multiplier_0_n_32_296));
  FA_X1_LVT multiplier_0_i_32_299 (.CO(multiplier_0_n_32_312), .S(
      multiplier_0_n_32_311), .A(multiplier_0_n_32_276), .B(
      multiplier_0_n_32_304), .CI(multiplier_0_n_32_297));
  FA_X1_LVT multiplier_0_i_32_326 (.CO(multiplier_0_n_32_344), .S(
      multiplier_0_n_32_343), .A(multiplier_0_n_32_318), .B(
      multiplier_0_n_32_339), .CI(multiplier_0_n_32_312));
  FA_X1_LVT multiplier_0_i_32_353 (.CO(multiplier_0_n_32_376), .S(
      multiplier_0_n_32_375), .A(multiplier_0_n_32_344), .B(
      multiplier_0_n_32_371), .CI(multiplier_0_n_32_373));
  XNOR2_X1_LVT multiplier_0_i_32_276 (.ZN(multiplier_0_n_32_287), .A(
      multiplier_0_n_32_137), .B(multiplier_0_n_32_121));
  XNOR2_X1_LVT multiplier_0_i_32_277 (.ZN(multiplier_0_n_32_288), .A(
      multiplier_0_n_32_287), .B(multiplier_0_n_32_105));
  OR2_X1_LVT multiplier_0_i_32_239 (.ZN(multiplier_0_n_32_244), .A1(
      multiplier_0_n_32_7), .A2(multiplier_0_n_32_23));
  INV_X1_LVT multiplier_0_i_32_241 (.ZN(multiplier_0_n_32_246), .A(
      multiplier_0_n_32_23));
  NAND2_X1_LVT multiplier_0_i_32_240 (.ZN(multiplier_0_n_32_245), .A1(
      multiplier_0_n_32_211), .A2(multiplier_0_n_32_246));
  INV_X1_LVT multiplier_0_i_32_243 (.ZN(multiplier_0_n_32_248), .A(
      multiplier_0_n_32_7));
  NAND2_X1_LVT multiplier_0_i_32_242 (.ZN(multiplier_0_n_32_247), .A1(
      multiplier_0_n_32_211), .A2(multiplier_0_n_32_248));
  NAND3_X1_LVT multiplier_0_i_32_238 (.ZN(multiplier_0_n_32_243), .A1(
      multiplier_0_n_32_244), .A2(multiplier_0_n_32_245), .A3(
      multiplier_0_n_32_247));
  XNOR2_X1_LVT multiplier_0_i_32_258 (.ZN(multiplier_0_n_32_266), .A(
      multiplier_0_n_32_56), .B(multiplier_0_n_32_40));
  XNOR2_X1_LVT multiplier_0_i_32_259 (.ZN(multiplier_0_n_32_267), .A(
      multiplier_0_n_32_266), .B(multiplier_0_n_32_24));
  INV_X1_LVT multiplier_0_i_32_260 (.ZN(multiplier_0_n_32_268), .A(
      multiplier_0_n_32_267));
  XNOR2_X1_LVT multiplier_0_i_32_251 (.ZN(multiplier_0_n_32_259), .A(
      multiplier_0_n_32_104), .B(multiplier_0_n_32_88));
  XNOR2_X1_LVT multiplier_0_i_32_252 (.ZN(multiplier_0_n_32_260), .A(
      multiplier_0_n_32_259), .B(multiplier_0_n_32_72));
  INV_X1_LVT multiplier_0_i_32_253 (.ZN(multiplier_0_n_32_261), .A(
      multiplier_0_n_32_260));
  FA_X1_LVT multiplier_0_i_32_273 (.CO(multiplier_0_n_32_282), .S(
      multiplier_0_n_32_281), .A(multiplier_0_n_32_243), .B(
      multiplier_0_n_32_268), .CI(multiplier_0_n_32_261));
  FA_X1_LVT multiplier_0_i_32_300 (.CO(multiplier_0_n_32_314), .S(
      multiplier_0_n_32_313), .A(multiplier_0_n_32_288), .B(
      multiplier_0_n_32_309), .CI(multiplier_0_n_32_282));
  FA_X1_LVT multiplier_0_i_32_327 (.CO(multiplier_0_n_32_346), .S(
      multiplier_0_n_32_345), .A(multiplier_0_n_32_314), .B(
      multiplier_0_n_32_341), .CI(multiplier_0_n_32_343));
  XNOR2_X1_LVT multiplier_0_i_32_247 (.ZN(multiplier_0_n_32_255), .A(
      multiplier_0_n_32_136), .B(multiplier_0_n_32_120));
  INV_X1_LVT multiplier_0_i_32_248 (.ZN(multiplier_0_n_32_256), .A(
      multiplier_0_n_32_255));
  XNOR2_X1_LVT multiplier_0_i_32_265 (.ZN(multiplier_0_n_32_273), .A(
      multiplier_0_n_32_8), .B(multiplier_0_n_32_237));
  XNOR2_X1_LVT multiplier_0_i_32_266 (.ZN(multiplier_0_n_32_274), .A(
      multiplier_0_n_32_273), .B(multiplier_0_n_32_230));
  INV_X1_LVT multiplier_0_i_32_267 (.ZN(multiplier_0_n_32_275), .A(
      multiplier_0_n_32_274));
  FA_X1_LVT multiplier_0_i_32_274 (.CO(multiplier_0_n_32_284), .S(
      multiplier_0_n_32_283), .A(multiplier_0_n_32_256), .B(
      multiplier_0_n_32_275), .CI(multiplier_0_n_32_250));
  FA_X1_LVT multiplier_0_i_32_301 (.CO(multiplier_0_n_32_316), .S(
      multiplier_0_n_32_315), .A(multiplier_0_n_32_284), .B(
      multiplier_0_n_32_311), .CI(multiplier_0_n_32_313));
  FA_X1_LVT multiplier_0_i_32_275 (.CO(multiplier_0_n_32_286), .S(
      multiplier_0_n_32_285), .A(multiplier_0_n_32_254), .B(
      multiplier_0_n_32_252), .CI(multiplier_0_n_32_281));
  FA_X1_LVT multiplier_0_i_32_602 (.CO(multiplier_0_n_32_659), .S(
      multiplier_0_n_50), .A(multiplier_0_n_32_283), .B(multiplier_0_n_32_285), 
      .CI(multiplier_0_n_32_658));
  FA_X1_LVT multiplier_0_i_32_603 (.CO(multiplier_0_n_32_660), .S(
      multiplier_0_n_51), .A(multiplier_0_n_32_286), .B(multiplier_0_n_32_315), 
      .CI(multiplier_0_n_32_659));
  FA_X1_LVT multiplier_0_i_32_604 (.CO(multiplier_0_n_32_661), .S(
      multiplier_0_n_52), .A(multiplier_0_n_32_316), .B(multiplier_0_n_32_345), 
      .CI(multiplier_0_n_32_660));
  FA_X1_LVT multiplier_0_i_32_605 (.CO(multiplier_0_n_32_662), .S(
      multiplier_0_n_53), .A(multiplier_0_n_32_346), .B(multiplier_0_n_32_375), 
      .CI(multiplier_0_n_32_661));
  FA_X1_LVT multiplier_0_i_32_606 (.CO(multiplier_0_n_32_663), .S(
      multiplier_0_n_54), .A(multiplier_0_n_32_376), .B(multiplier_0_n_32_405), 
      .CI(multiplier_0_n_32_662));
  FA_X1_LVT multiplier_0_i_32_607 (.CO(multiplier_0_n_32_664), .S(
      multiplier_0_n_55), .A(multiplier_0_n_32_406), .B(multiplier_0_n_32_435), 
      .CI(multiplier_0_n_32_663));
  FA_X1_LVT multiplier_0_i_32_608 (.CO(multiplier_0_n_32_665), .S(
      multiplier_0_n_56), .A(multiplier_0_n_32_436), .B(multiplier_0_n_32_465), 
      .CI(multiplier_0_n_32_664));
  FA_X1_LVT multiplier_0_i_32_609 (.CO(multiplier_0_n_32_666), .S(
      multiplier_0_n_57), .A(multiplier_0_n_32_466), .B(multiplier_0_n_32_495), 
      .CI(multiplier_0_n_32_665));
  INV_X1_LVT multiplier_0_i_34_31 (.ZN(multiplier_0_n_34_16), .A(
      multiplier_0_n_57));
  OAI22_X1_LVT multiplier_0_i_34_32 (.ZN(multiplier_0_product_xp[15]), .A1(
      multiplier_0_n_34_8), .A2(multiplier_0_n_34_7), .B1(multiplier_0_n_34_16), 
      .B2(multiplier_0_cycle[0]));
  INV_X1_LVT multiplier_0_i_34_12 (.ZN(multiplier_0_n_34_6), .A(
      multiplier_0_n_48));
  INV_X1_LVT multiplier_0_i_34_29 (.ZN(multiplier_0_n_34_15), .A(
      multiplier_0_n_56));
  OAI22_X1_LVT multiplier_0_i_34_30 (.ZN(multiplier_0_product_xp[14]), .A1(
      multiplier_0_n_34_8), .A2(multiplier_0_n_34_6), .B1(multiplier_0_n_34_15), 
      .B2(multiplier_0_cycle[0]));
  AOI22_X1_LVT multiplier_0_i_45_29 (.ZN(multiplier_0_n_45_15), .A1(
      multiplier_0_n_45_0), .A2(multiplier_0_n_136), .B1(multiplier_0_reslo_wr), 
      .B2(multiplier_0_per_din_msk[14]));
  INV_X1_LVT multiplier_0_i_45_30 (.ZN(multiplier_0_n_119), .A(
      multiplier_0_n_45_15));
  OR2_X1_LVT multiplier_0_i_23_0 (.ZN(multiplier_0_result_wr), .A1(
      multiplier_0_cycle[0]), .A2(multiplier_0_cycle[1]));
  INV_X1_LVT multiplier_0_i_39_1 (.ZN(multiplier_0_n_39_1), .A(
      multiplier_0_result_wr));
  INV_X1_LVT multiplier_0_i_39_0 (.ZN(multiplier_0_n_39_0), .A(
      multiplier_0_result_clr));
  NAND2_X1_LVT multiplier_0_i_39_2 (.ZN(multiplier_0_n_69), .A1(
      multiplier_0_n_39_1), .A2(multiplier_0_n_39_0));
  INV_X1_LVT multiplier_0_i_46_1 (.ZN(multiplier_0_n_46_1), .A(multiplier_0_n_69));
  INV_X1_LVT multiplier_0_i_46_0 (.ZN(multiplier_0_n_46_0), .A(
      multiplier_0_reslo_wr));
  NAND2_X1_LVT multiplier_0_i_46_2 (.ZN(multiplier_0_n_121), .A1(
      multiplier_0_n_46_1), .A2(multiplier_0_n_46_0));
  CLKGATETST_X1_LVT multiplier_0_clk_gate_reslo_reg (.GCK(multiplier_0_n_88), 
      .CK(mclk), .E(multiplier_0_n_121), .SE(1'b0));
  DFFR_X1_LVT \multiplier_0_reslo_reg[14] (.Q(multiplier_0_n_90), .QN(), .CK(
      multiplier_0_n_88), .D(multiplier_0_n_119), .RN(multiplier_0_n_38));
  INV_X1_LVT multiplier_0_i_34_10 (.ZN(multiplier_0_n_34_5), .A(
      multiplier_0_n_47));
  INV_X1_LVT multiplier_0_i_34_27 (.ZN(multiplier_0_n_34_14), .A(
      multiplier_0_n_55));
  OAI22_X1_LVT multiplier_0_i_34_28 (.ZN(multiplier_0_product_xp[13]), .A1(
      multiplier_0_n_34_8), .A2(multiplier_0_n_34_5), .B1(multiplier_0_n_34_14), 
      .B2(multiplier_0_cycle[0]));
  AOI22_X1_LVT multiplier_0_i_45_27 (.ZN(multiplier_0_n_45_14), .A1(
      multiplier_0_n_45_0), .A2(multiplier_0_n_135), .B1(multiplier_0_reslo_wr), 
      .B2(multiplier_0_per_din_msk[13]));
  INV_X1_LVT multiplier_0_i_45_28 (.ZN(multiplier_0_n_118), .A(
      multiplier_0_n_45_14));
  DFFR_X1_LVT \multiplier_0_reslo_reg[13] (.Q(multiplier_0_n_91), .QN(), .CK(
      multiplier_0_n_88), .D(multiplier_0_n_118), .RN(multiplier_0_n_38));
  INV_X1_LVT multiplier_0_i_34_8 (.ZN(multiplier_0_n_34_4), .A(multiplier_0_n_46));
  INV_X1_LVT multiplier_0_i_34_25 (.ZN(multiplier_0_n_34_13), .A(
      multiplier_0_n_54));
  OAI22_X1_LVT multiplier_0_i_34_26 (.ZN(multiplier_0_product_xp[12]), .A1(
      multiplier_0_n_34_8), .A2(multiplier_0_n_34_4), .B1(multiplier_0_n_34_13), 
      .B2(multiplier_0_cycle[0]));
  AOI22_X1_LVT multiplier_0_i_45_25 (.ZN(multiplier_0_n_45_13), .A1(
      multiplier_0_n_45_0), .A2(multiplier_0_n_134), .B1(multiplier_0_reslo_wr), 
      .B2(multiplier_0_per_din_msk[12]));
  INV_X1_LVT multiplier_0_i_45_26 (.ZN(multiplier_0_n_117), .A(
      multiplier_0_n_45_13));
  DFFR_X1_LVT \multiplier_0_reslo_reg[12] (.Q(multiplier_0_n_92), .QN(), .CK(
      multiplier_0_n_88), .D(multiplier_0_n_117), .RN(multiplier_0_n_38));
  INV_X1_LVT multiplier_0_i_34_6 (.ZN(multiplier_0_n_34_3), .A(multiplier_0_n_45));
  INV_X1_LVT multiplier_0_i_34_23 (.ZN(multiplier_0_n_34_12), .A(
      multiplier_0_n_53));
  OAI22_X1_LVT multiplier_0_i_34_24 (.ZN(multiplier_0_product_xp[11]), .A1(
      multiplier_0_n_34_8), .A2(multiplier_0_n_34_3), .B1(multiplier_0_n_34_12), 
      .B2(multiplier_0_cycle[0]));
  AOI22_X1_LVT multiplier_0_i_45_23 (.ZN(multiplier_0_n_45_12), .A1(
      multiplier_0_n_45_0), .A2(multiplier_0_n_133), .B1(multiplier_0_reslo_wr), 
      .B2(multiplier_0_per_din_msk[11]));
  INV_X1_LVT multiplier_0_i_45_24 (.ZN(multiplier_0_n_116), .A(
      multiplier_0_n_45_12));
  DFFR_X1_LVT \multiplier_0_reslo_reg[11] (.Q(multiplier_0_n_93), .QN(), .CK(
      multiplier_0_n_88), .D(multiplier_0_n_116), .RN(multiplier_0_n_38));
  XNOR2_X1_LVT multiplier_0_i_32_589 (.ZN(multiplier_0_n_32_647), .A(
      multiplier_0_n_32_2), .B(multiplier_0_n_32_153));
  XNOR2_X1_LVT multiplier_0_i_32_590 (.ZN(multiplier_0_n_32_648), .A(
      multiplier_0_n_32_647), .B(multiplier_0_n_32_646));
  INV_X1_LVT multiplier_0_i_32_591 (.ZN(multiplier_0_n_44), .A(
      multiplier_0_n_32_648));
  INV_X1_LVT multiplier_0_i_34_4 (.ZN(multiplier_0_n_34_2), .A(multiplier_0_n_44));
  INV_X1_LVT multiplier_0_i_34_21 (.ZN(multiplier_0_n_34_11), .A(
      multiplier_0_n_52));
  OAI22_X1_LVT multiplier_0_i_34_22 (.ZN(multiplier_0_product_xp[10]), .A1(
      multiplier_0_n_34_8), .A2(multiplier_0_n_34_2), .B1(multiplier_0_n_34_11), 
      .B2(multiplier_0_cycle[0]));
  AOI22_X1_LVT multiplier_0_i_45_21 (.ZN(multiplier_0_n_45_11), .A1(
      multiplier_0_n_45_0), .A2(multiplier_0_n_132), .B1(multiplier_0_reslo_wr), 
      .B2(multiplier_0_per_din_msk[10]));
  INV_X1_LVT multiplier_0_i_45_22 (.ZN(multiplier_0_n_115), .A(
      multiplier_0_n_45_11));
  DFFR_X1_LVT \multiplier_0_reslo_reg[10] (.Q(multiplier_0_n_94), .QN(), .CK(
      multiplier_0_n_88), .D(multiplier_0_n_115), .RN(multiplier_0_n_38));
  XNOR2_X1_LVT multiplier_0_i_32_586 (.ZN(multiplier_0_n_32_645), .A(
      multiplier_0_n_32_17), .B(multiplier_0_n_32_1));
  INV_X1_LVT multiplier_0_i_32_587 (.ZN(multiplier_0_n_43), .A(
      multiplier_0_n_32_645));
  INV_X1_LVT multiplier_0_i_34_2 (.ZN(multiplier_0_n_34_1), .A(multiplier_0_n_43));
  INV_X1_LVT multiplier_0_i_34_19 (.ZN(multiplier_0_n_34_10), .A(
      multiplier_0_n_51));
  OAI22_X1_LVT multiplier_0_i_34_20 (.ZN(multiplier_0_product_xp[9]), .A1(
      multiplier_0_n_34_8), .A2(multiplier_0_n_34_1), .B1(multiplier_0_n_34_10), 
      .B2(multiplier_0_cycle[0]));
  AOI22_X1_LVT multiplier_0_i_45_19 (.ZN(multiplier_0_n_45_10), .A1(
      multiplier_0_n_45_0), .A2(multiplier_0_n_131), .B1(multiplier_0_reslo_wr), 
      .B2(multiplier_0_per_din_msk[9]));
  INV_X1_LVT multiplier_0_i_45_20 (.ZN(multiplier_0_n_114), .A(
      multiplier_0_n_45_10));
  DFFR_X1_LVT \multiplier_0_reslo_reg[9] (.Q(multiplier_0_n_95), .QN(), .CK(
      multiplier_0_n_88), .D(multiplier_0_n_114), .RN(multiplier_0_n_38));
  NAND2_X1_LVT multiplier_0_i_32_0 (.ZN(multiplier_0_n_32_0), .A1(
      multiplier_0_op2_xp[0]), .A2(multiplier_0_op1[0]));
  INV_X1_LVT multiplier_0_i_32_585 (.ZN(multiplier_0_n_42), .A(
      multiplier_0_n_32_0));
  INV_X1_LVT multiplier_0_i_34_0 (.ZN(multiplier_0_n_34_0), .A(multiplier_0_n_42));
  INV_X1_LVT multiplier_0_i_34_17 (.ZN(multiplier_0_n_34_9), .A(
      multiplier_0_n_50));
  OAI22_X1_LVT multiplier_0_i_34_18 (.ZN(multiplier_0_product_xp[8]), .A1(
      multiplier_0_n_34_0), .A2(multiplier_0_n_34_8), .B1(multiplier_0_n_34_9), 
      .B2(multiplier_0_cycle[0]));
  AOI22_X1_LVT multiplier_0_i_45_17 (.ZN(multiplier_0_n_45_9), .A1(
      multiplier_0_n_45_0), .A2(multiplier_0_n_130), .B1(multiplier_0_reslo_wr), 
      .B2(multiplier_0_per_din_msk[8]));
  INV_X1_LVT multiplier_0_i_45_18 (.ZN(multiplier_0_n_113), .A(
      multiplier_0_n_45_9));
  DFFR_X1_LVT \multiplier_0_reslo_reg[8] (.Q(multiplier_0_n_96), .QN(), .CK(
      multiplier_0_n_88), .D(multiplier_0_n_113), .RN(multiplier_0_n_38));
  NOR2_X1_LVT multiplier_0_i_34_15 (.ZN(multiplier_0_product_xp[7]), .A1(
      multiplier_0_n_34_7), .A2(multiplier_0_cycle[0]));
  AOI22_X1_LVT multiplier_0_i_45_15 (.ZN(multiplier_0_n_45_8), .A1(
      multiplier_0_n_45_0), .A2(multiplier_0_n_129), .B1(multiplier_0_reslo_wr), 
      .B2(per_din[7]));
  INV_X1_LVT multiplier_0_i_45_16 (.ZN(multiplier_0_n_112), .A(
      multiplier_0_n_45_8));
  DFFR_X1_LVT \multiplier_0_reslo_reg[7] (.Q(multiplier_0_n_97), .QN(), .CK(
      multiplier_0_n_88), .D(multiplier_0_n_112), .RN(multiplier_0_n_38));
  NOR2_X1_LVT multiplier_0_i_34_13 (.ZN(multiplier_0_product_xp[6]), .A1(
      multiplier_0_n_34_6), .A2(multiplier_0_cycle[0]));
  AOI22_X1_LVT multiplier_0_i_45_13 (.ZN(multiplier_0_n_45_7), .A1(
      multiplier_0_n_45_0), .A2(multiplier_0_n_128), .B1(multiplier_0_reslo_wr), 
      .B2(per_din[6]));
  INV_X1_LVT multiplier_0_i_45_14 (.ZN(multiplier_0_n_111), .A(
      multiplier_0_n_45_7));
  DFFR_X1_LVT \multiplier_0_reslo_reg[6] (.Q(multiplier_0_n_98), .QN(), .CK(
      multiplier_0_n_88), .D(multiplier_0_n_111), .RN(multiplier_0_n_38));
  NOR2_X1_LVT multiplier_0_i_34_11 (.ZN(multiplier_0_product_xp[5]), .A1(
      multiplier_0_n_34_5), .A2(multiplier_0_cycle[0]));
  AOI22_X1_LVT multiplier_0_i_45_11 (.ZN(multiplier_0_n_45_6), .A1(
      multiplier_0_n_45_0), .A2(multiplier_0_n_127), .B1(multiplier_0_reslo_wr), 
      .B2(per_din[5]));
  INV_X1_LVT multiplier_0_i_45_12 (.ZN(multiplier_0_n_110), .A(
      multiplier_0_n_45_6));
  DFFR_X1_LVT \multiplier_0_reslo_reg[5] (.Q(multiplier_0_n_99), .QN(), .CK(
      multiplier_0_n_88), .D(multiplier_0_n_110), .RN(multiplier_0_n_38));
  NOR2_X1_LVT multiplier_0_i_34_9 (.ZN(multiplier_0_product_xp[4]), .A1(
      multiplier_0_n_34_4), .A2(multiplier_0_cycle[0]));
  AOI22_X1_LVT multiplier_0_i_45_9 (.ZN(multiplier_0_n_45_5), .A1(
      multiplier_0_n_45_0), .A2(multiplier_0_n_126), .B1(multiplier_0_reslo_wr), 
      .B2(per_din[4]));
  INV_X1_LVT multiplier_0_i_45_10 (.ZN(multiplier_0_n_109), .A(
      multiplier_0_n_45_5));
  DFFR_X1_LVT \multiplier_0_reslo_reg[4] (.Q(multiplier_0_n_100), .QN(), .CK(
      multiplier_0_n_88), .D(multiplier_0_n_109), .RN(multiplier_0_n_38));
  NOR2_X1_LVT multiplier_0_i_34_7 (.ZN(multiplier_0_product_xp[3]), .A1(
      multiplier_0_n_34_3), .A2(multiplier_0_cycle[0]));
  AOI22_X1_LVT multiplier_0_i_45_7 (.ZN(multiplier_0_n_45_4), .A1(
      multiplier_0_n_45_0), .A2(multiplier_0_n_125), .B1(multiplier_0_reslo_wr), 
      .B2(per_din[3]));
  INV_X1_LVT multiplier_0_i_45_8 (.ZN(multiplier_0_n_108), .A(
      multiplier_0_n_45_4));
  DFFR_X1_LVT \multiplier_0_reslo_reg[3] (.Q(multiplier_0_n_101), .QN(), .CK(
      multiplier_0_n_88), .D(multiplier_0_n_108), .RN(multiplier_0_n_38));
  NOR2_X1_LVT multiplier_0_i_34_5 (.ZN(multiplier_0_product_xp[2]), .A1(
      multiplier_0_n_34_2), .A2(multiplier_0_cycle[0]));
  AOI22_X1_LVT multiplier_0_i_45_5 (.ZN(multiplier_0_n_45_3), .A1(
      multiplier_0_n_45_0), .A2(multiplier_0_n_124), .B1(multiplier_0_reslo_wr), 
      .B2(per_din[2]));
  INV_X1_LVT multiplier_0_i_45_6 (.ZN(multiplier_0_n_107), .A(
      multiplier_0_n_45_3));
  DFFR_X1_LVT \multiplier_0_reslo_reg[2] (.Q(multiplier_0_n_102), .QN(), .CK(
      multiplier_0_n_88), .D(multiplier_0_n_107), .RN(multiplier_0_n_38));
  NOR2_X1_LVT multiplier_0_i_34_3 (.ZN(multiplier_0_product_xp[1]), .A1(
      multiplier_0_n_34_1), .A2(multiplier_0_cycle[0]));
  AOI22_X1_LVT multiplier_0_i_45_3 (.ZN(multiplier_0_n_45_2), .A1(
      multiplier_0_n_45_0), .A2(multiplier_0_n_123), .B1(multiplier_0_reslo_wr), 
      .B2(per_din[1]));
  INV_X1_LVT multiplier_0_i_45_4 (.ZN(multiplier_0_n_106), .A(
      multiplier_0_n_45_2));
  DFFR_X1_LVT \multiplier_0_reslo_reg[1] (.Q(multiplier_0_n_103), .QN(), .CK(
      multiplier_0_n_88), .D(multiplier_0_n_106), .RN(multiplier_0_n_38));
  NOR2_X1_LVT multiplier_0_i_34_1 (.ZN(multiplier_0_product_xp[0]), .A1(
      multiplier_0_n_34_0), .A2(multiplier_0_cycle[0]));
  AOI22_X1_LVT multiplier_0_i_45_1 (.ZN(multiplier_0_n_45_1), .A1(
      multiplier_0_n_45_0), .A2(multiplier_0_n_122), .B1(per_din[0]), .B2(
      multiplier_0_reslo_wr));
  INV_X1_LVT multiplier_0_i_45_2 (.ZN(multiplier_0_n_105), .A(
      multiplier_0_n_45_1));
  DFFR_X1_LVT \multiplier_0_reslo_reg[0] (.Q(multiplier_0_n_104), .QN(), .CK(
      multiplier_0_n_88), .D(multiplier_0_n_105), .RN(multiplier_0_n_38));
  HA_X1_LVT multiplier_0_i_48_0 (.CO(multiplier_0_n_48_0), .S(multiplier_0_n_122), 
      .A(multiplier_0_product_xp[0]), .B(multiplier_0_n_104));
  FA_X1_LVT multiplier_0_i_48_1 (.CO(multiplier_0_n_48_1), .S(multiplier_0_n_123), 
      .A(multiplier_0_product_xp[1]), .B(multiplier_0_n_103), .CI(
      multiplier_0_n_48_0));
  FA_X1_LVT multiplier_0_i_48_2 (.CO(multiplier_0_n_48_2), .S(multiplier_0_n_124), 
      .A(multiplier_0_product_xp[2]), .B(multiplier_0_n_102), .CI(
      multiplier_0_n_48_1));
  FA_X1_LVT multiplier_0_i_48_3 (.CO(multiplier_0_n_48_3), .S(multiplier_0_n_125), 
      .A(multiplier_0_product_xp[3]), .B(multiplier_0_n_101), .CI(
      multiplier_0_n_48_2));
  FA_X1_LVT multiplier_0_i_48_4 (.CO(multiplier_0_n_48_4), .S(multiplier_0_n_126), 
      .A(multiplier_0_product_xp[4]), .B(multiplier_0_n_100), .CI(
      multiplier_0_n_48_3));
  FA_X1_LVT multiplier_0_i_48_5 (.CO(multiplier_0_n_48_5), .S(multiplier_0_n_127), 
      .A(multiplier_0_product_xp[5]), .B(multiplier_0_n_99), .CI(
      multiplier_0_n_48_4));
  FA_X1_LVT multiplier_0_i_48_6 (.CO(multiplier_0_n_48_6), .S(multiplier_0_n_128), 
      .A(multiplier_0_product_xp[6]), .B(multiplier_0_n_98), .CI(
      multiplier_0_n_48_5));
  FA_X1_LVT multiplier_0_i_48_7 (.CO(multiplier_0_n_48_7), .S(multiplier_0_n_129), 
      .A(multiplier_0_product_xp[7]), .B(multiplier_0_n_97), .CI(
      multiplier_0_n_48_6));
  FA_X1_LVT multiplier_0_i_48_8 (.CO(multiplier_0_n_48_8), .S(multiplier_0_n_130), 
      .A(multiplier_0_product_xp[8]), .B(multiplier_0_n_96), .CI(
      multiplier_0_n_48_7));
  FA_X1_LVT multiplier_0_i_48_9 (.CO(multiplier_0_n_48_9), .S(multiplier_0_n_131), 
      .A(multiplier_0_product_xp[9]), .B(multiplier_0_n_95), .CI(
      multiplier_0_n_48_8));
  FA_X1_LVT multiplier_0_i_48_10 (.CO(multiplier_0_n_48_10), .S(
      multiplier_0_n_132), .A(multiplier_0_product_xp[10]), .B(multiplier_0_n_94), 
      .CI(multiplier_0_n_48_9));
  FA_X1_LVT multiplier_0_i_48_11 (.CO(multiplier_0_n_48_11), .S(
      multiplier_0_n_133), .A(multiplier_0_product_xp[11]), .B(multiplier_0_n_93), 
      .CI(multiplier_0_n_48_10));
  FA_X1_LVT multiplier_0_i_48_12 (.CO(multiplier_0_n_48_12), .S(
      multiplier_0_n_134), .A(multiplier_0_product_xp[12]), .B(multiplier_0_n_92), 
      .CI(multiplier_0_n_48_11));
  FA_X1_LVT multiplier_0_i_48_13 (.CO(multiplier_0_n_48_13), .S(
      multiplier_0_n_135), .A(multiplier_0_product_xp[13]), .B(multiplier_0_n_91), 
      .CI(multiplier_0_n_48_12));
  FA_X1_LVT multiplier_0_i_48_14 (.CO(multiplier_0_n_48_14), .S(
      multiplier_0_n_136), .A(multiplier_0_product_xp[14]), .B(multiplier_0_n_90), 
      .CI(multiplier_0_n_48_13));
  FA_X1_LVT multiplier_0_i_48_15 (.CO(multiplier_0_n_48_15), .S(
      multiplier_0_n_137), .A(multiplier_0_product_xp[15]), .B(multiplier_0_n_89), 
      .CI(multiplier_0_n_48_14));
  AOI22_X1_LVT multiplier_0_i_45_31 (.ZN(multiplier_0_n_45_16), .A1(
      multiplier_0_n_45_0), .A2(multiplier_0_n_137), .B1(multiplier_0_reslo_wr), 
      .B2(multiplier_0_per_din_msk[15]));
  INV_X1_LVT multiplier_0_i_45_32 (.ZN(multiplier_0_n_120), .A(
      multiplier_0_n_45_16));
  DFFR_X1_LVT \multiplier_0_reslo_reg[15] (.Q(multiplier_0_n_89), .QN(), .CK(
      multiplier_0_n_88), .D(multiplier_0_n_120), .RN(multiplier_0_n_38));
  AOI22_X1_LVT multiplier_0_i_60_93 (.ZN(multiplier_0_n_60_78), .A1(
      multiplier_0_n_60_0), .A2(multiplier_0_n_89), .B1(multiplier_0_cycle[1]), 
      .B2(multiplier_0_n_137));
  NOR2_X1_LVT multiplier_0_i_1_0 (.ZN(multiplier_0_n_0), .A1(per_we[0]), .A2(
      per_we[1]));
  AND2_X1_LVT multiplier_0_i_2_0 (.ZN(multiplier_0_reg_read), .A1(
      multiplier_0_n_0), .A2(multiplier_0_reg_sel));
  AND2_X1_LVT multiplier_0_i_4_5 (.ZN(multiplier_0_n_13), .A1(
      multiplier_0_reg_read), .A2(multiplier_0_n_6));
  INV_X1_LVT multiplier_0_i_60_2 (.ZN(multiplier_0_n_60_2), .A(multiplier_0_n_13));
  NOR2_X1_LVT multiplier_0_i_60_94 (.ZN(multiplier_0_n_60_79), .A1(
      multiplier_0_n_60_78), .A2(multiplier_0_n_60_2));
  AND2_X1_LVT multiplier_0_i_4_0 (.ZN(multiplier_0_n_9), .A1(multiplier_0_n_1), 
      .A2(multiplier_0_reg_read));
  AND2_X1_LVT multiplier_0_i_4_3 (.ZN(multiplier_0_n_11), .A1(
      multiplier_0_reg_read), .A2(multiplier_0_n_4));
  AND2_X1_LVT multiplier_0_i_4_2 (.ZN(multiplier_0_reg_rd1), .A1(
      multiplier_0_reg_read), .A2(multiplier_0_n_3));
  AND2_X1_LVT multiplier_0_i_4_1 (.ZN(multiplier_0_n_10), .A1(
      multiplier_0_reg_read), .A2(multiplier_0_n_2));
  OR4_X1_LVT multiplier_0_i_59_0 (.ZN(multiplier_0_n_150), .A1(multiplier_0_n_9), 
      .A2(multiplier_0_n_11), .A3(multiplier_0_reg_rd1), .A4(multiplier_0_n_10));
  AND2_X1_LVT multiplier_0_i_60_95 (.ZN(multiplier_0_n_60_80), .A1(
      multiplier_0_n_150), .A2(multiplier_0_op1[15]));
  INV_X1_LVT multiplier_0_i_57_0 (.ZN(multiplier_0_n_57_0), .A(
      multiplier_0_cycle[1]));
  INV_X1_LVT multiplier_0_i_52_0 (.ZN(multiplier_0_n_52_0), .A(
      multiplier_0_op2_wr));
  NAND2_X1_LVT multiplier_0_i_32_151 (.ZN(multiplier_0_n_32_151), .A1(
      multiplier_0_op2_xp[8]), .A2(multiplier_0_op1[15]));
  AND2_X1_LVT multiplier_0_i_31_0 (.ZN(multiplier_0_op1_xp[16]), .A1(
      multiplier_0_op1[15]), .A2(multiplier_0_sign_sel));
  NAND2_X1_LVT multiplier_0_i_32_135 (.ZN(multiplier_0_n_32_135), .A1(
      multiplier_0_op2_xp[7]), .A2(multiplier_0_op1_xp[16]));
  XNOR2_X1_LVT multiplier_0_i_32_583 (.ZN(multiplier_0_n_32_643), .A(
      multiplier_0_n_32_151), .B(multiplier_0_n_32_135));
  NAND2_X1_LVT multiplier_0_i_32_150 (.ZN(multiplier_0_n_32_150), .A1(
      multiplier_0_op2_xp[8]), .A2(multiplier_0_op1[14]));
  NAND2_X1_LVT multiplier_0_i_32_134 (.ZN(multiplier_0_n_32_134), .A1(
      multiplier_0_op2_xp[7]), .A2(multiplier_0_op1[15]));
  INV_X1_LVT multiplier_0_i_32_579 (.ZN(multiplier_0_n_32_638), .A(
      multiplier_0_n_32_134));
  NAND2_X1_LVT multiplier_0_i_32_578 (.ZN(multiplier_0_n_32_637), .A1(
      multiplier_0_n_32_150), .A2(multiplier_0_n_32_638));
  NAND2_X1_LVT multiplier_0_i_32_118 (.ZN(multiplier_0_n_32_118), .A1(
      multiplier_0_op2_xp[6]), .A2(multiplier_0_op1_xp[16]));
  NAND2_X1_LVT multiplier_0_i_32_580 (.ZN(multiplier_0_n_32_639), .A1(
      multiplier_0_n_32_118), .A2(multiplier_0_n_32_150));
  NAND2_X1_LVT multiplier_0_i_32_581 (.ZN(multiplier_0_n_32_640), .A1(
      multiplier_0_n_32_118), .A2(multiplier_0_n_32_638));
  NAND3_X1_LVT multiplier_0_i_32_577 (.ZN(multiplier_0_n_32_636), .A1(
      multiplier_0_n_32_637), .A2(multiplier_0_n_32_639), .A3(
      multiplier_0_n_32_640));
  XNOR2_X1_LVT multiplier_0_i_32_584 (.ZN(multiplier_0_n_32_644), .A(
      multiplier_0_n_32_643), .B(multiplier_0_n_32_636));
  NAND2_X1_LVT multiplier_0_i_32_149 (.ZN(multiplier_0_n_32_149), .A1(
      multiplier_0_op2_xp[8]), .A2(multiplier_0_op1[13]));
  NAND2_X1_LVT multiplier_0_i_32_133 (.ZN(multiplier_0_n_32_133), .A1(
      multiplier_0_op2_xp[7]), .A2(multiplier_0_op1[14]));
  INV_X1_LVT multiplier_0_i_32_568 (.ZN(multiplier_0_n_32_625), .A(
      multiplier_0_n_32_133));
  NAND2_X1_LVT multiplier_0_i_32_567 (.ZN(multiplier_0_n_32_624), .A1(
      multiplier_0_n_32_149), .A2(multiplier_0_n_32_625));
  NAND2_X1_LVT multiplier_0_i_32_117 (.ZN(multiplier_0_n_32_117), .A1(
      multiplier_0_op2_xp[6]), .A2(multiplier_0_op1[15]));
  INV_X1_LVT multiplier_0_i_32_570 (.ZN(multiplier_0_n_32_627), .A(
      multiplier_0_n_32_117));
  NAND2_X1_LVT multiplier_0_i_32_569 (.ZN(multiplier_0_n_32_626), .A1(
      multiplier_0_n_32_149), .A2(multiplier_0_n_32_627));
  OR2_X1_LVT multiplier_0_i_32_571 (.ZN(multiplier_0_n_32_628), .A1(
      multiplier_0_n_32_117), .A2(multiplier_0_n_32_133));
  NAND3_X1_LVT multiplier_0_i_32_566 (.ZN(multiplier_0_n_32_623), .A1(
      multiplier_0_n_32_624), .A2(multiplier_0_n_32_626), .A3(
      multiplier_0_n_32_628));
  NAND2_X1_LVT multiplier_0_i_32_101 (.ZN(multiplier_0_n_32_101), .A1(
      multiplier_0_op2_xp[5]), .A2(multiplier_0_op1_xp[16]));
  NAND2_X1_LVT multiplier_0_i_32_148 (.ZN(multiplier_0_n_32_148), .A1(
      multiplier_0_op2_xp[8]), .A2(multiplier_0_op1[12]));
  NAND2_X1_LVT multiplier_0_i_32_132 (.ZN(multiplier_0_n_32_132), .A1(
      multiplier_0_op2_xp[7]), .A2(multiplier_0_op1[13]));
  INV_X1_LVT multiplier_0_i_32_550 (.ZN(multiplier_0_n_32_605), .A(
      multiplier_0_n_32_132));
  NAND2_X1_LVT multiplier_0_i_32_549 (.ZN(multiplier_0_n_32_604), .A1(
      multiplier_0_n_32_148), .A2(multiplier_0_n_32_605));
  NAND2_X1_LVT multiplier_0_i_32_116 (.ZN(multiplier_0_n_32_116), .A1(
      multiplier_0_op2_xp[6]), .A2(multiplier_0_op1[14]));
  INV_X1_LVT multiplier_0_i_32_552 (.ZN(multiplier_0_n_32_607), .A(
      multiplier_0_n_32_116));
  NAND2_X1_LVT multiplier_0_i_32_551 (.ZN(multiplier_0_n_32_606), .A1(
      multiplier_0_n_32_148), .A2(multiplier_0_n_32_607));
  OR2_X1_LVT multiplier_0_i_32_553 (.ZN(multiplier_0_n_32_608), .A1(
      multiplier_0_n_32_116), .A2(multiplier_0_n_32_132));
  NAND3_X1_LVT multiplier_0_i_32_548 (.ZN(multiplier_0_n_32_603), .A1(
      multiplier_0_n_32_604), .A2(multiplier_0_n_32_606), .A3(
      multiplier_0_n_32_608));
  NAND2_X1_LVT multiplier_0_i_32_84 (.ZN(multiplier_0_n_32_84), .A1(
      multiplier_0_op2_xp[4]), .A2(multiplier_0_op1_xp[16]));
  NAND2_X1_LVT multiplier_0_i_32_100 (.ZN(multiplier_0_n_32_100), .A1(
      multiplier_0_op2_xp[5]), .A2(multiplier_0_op1[15]));
  INV_X1_LVT multiplier_0_i_32_559 (.ZN(multiplier_0_n_32_614), .A(
      multiplier_0_n_32_100));
  NAND2_X1_LVT multiplier_0_i_32_558 (.ZN(multiplier_0_n_32_613), .A1(
      multiplier_0_n_32_84), .A2(multiplier_0_n_32_614));
  NAND2_X1_LVT multiplier_0_i_32_83 (.ZN(multiplier_0_n_32_83), .A1(
      multiplier_0_op2_xp[4]), .A2(multiplier_0_op1[15]));
  NAND2_X1_LVT multiplier_0_i_32_99 (.ZN(multiplier_0_n_32_99), .A1(
      multiplier_0_op2_xp[5]), .A2(multiplier_0_op1[14]));
  OR2_X1_LVT multiplier_0_i_32_538 (.ZN(multiplier_0_n_32_590), .A1(
      multiplier_0_n_32_83), .A2(multiplier_0_n_32_99));
  NAND2_X1_LVT multiplier_0_i_32_67 (.ZN(multiplier_0_n_32_67), .A1(
      multiplier_0_op2_xp[3]), .A2(multiplier_0_op1_xp[16]));
  INV_X1_LVT multiplier_0_i_32_540 (.ZN(multiplier_0_n_32_592), .A(
      multiplier_0_n_32_99));
  NAND2_X1_LVT multiplier_0_i_32_539 (.ZN(multiplier_0_n_32_591), .A1(
      multiplier_0_n_32_67), .A2(multiplier_0_n_32_592));
  INV_X1_LVT multiplier_0_i_32_542 (.ZN(multiplier_0_n_32_594), .A(
      multiplier_0_n_32_83));
  NAND2_X1_LVT multiplier_0_i_32_541 (.ZN(multiplier_0_n_32_593), .A1(
      multiplier_0_n_32_67), .A2(multiplier_0_n_32_594));
  NAND3_X1_LVT multiplier_0_i_32_537 (.ZN(multiplier_0_n_32_589), .A1(
      multiplier_0_n_32_590), .A2(multiplier_0_n_32_591), .A3(
      multiplier_0_n_32_593));
  NAND2_X1_LVT multiplier_0_i_32_560 (.ZN(multiplier_0_n_32_615), .A1(
      multiplier_0_n_32_589), .A2(multiplier_0_n_32_614));
  NAND2_X1_LVT multiplier_0_i_32_561 (.ZN(multiplier_0_n_32_616), .A1(
      multiplier_0_n_32_589), .A2(multiplier_0_n_32_84));
  NAND3_X1_LVT multiplier_0_i_32_557 (.ZN(multiplier_0_n_32_612), .A1(
      multiplier_0_n_32_613), .A2(multiplier_0_n_32_615), .A3(
      multiplier_0_n_32_616));
  FA_X1_LVT multiplier_0_i_32_572 (.CO(multiplier_0_n_32_630), .S(
      multiplier_0_n_32_629), .A(multiplier_0_n_32_101), .B(
      multiplier_0_n_32_603), .CI(multiplier_0_n_32_612));
  XNOR2_X1_LVT multiplier_0_i_32_574 (.ZN(multiplier_0_n_32_633), .A(
      multiplier_0_n_32_150), .B(multiplier_0_n_32_134));
  XNOR2_X1_LVT multiplier_0_i_32_575 (.ZN(multiplier_0_n_32_634), .A(
      multiplier_0_n_32_633), .B(multiplier_0_n_32_118));
  INV_X1_LVT multiplier_0_i_32_576 (.ZN(multiplier_0_n_32_635), .A(
      multiplier_0_n_32_634));
  FA_X1_LVT multiplier_0_i_32_582 (.CO(multiplier_0_n_32_642), .S(
      multiplier_0_n_32_641), .A(multiplier_0_n_32_623), .B(
      multiplier_0_n_32_630), .CI(multiplier_0_n_32_635));
  XNOR2_X1_LVT multiplier_0_i_32_617 (.ZN(multiplier_0_n_32_674), .A(
      multiplier_0_n_32_644), .B(multiplier_0_n_32_642));
  XNOR2_X1_LVT multiplier_0_i_32_564 (.ZN(multiplier_0_n_32_621), .A(
      multiplier_0_n_32_149), .B(multiplier_0_n_32_133));
  XNOR2_X1_LVT multiplier_0_i_32_565 (.ZN(multiplier_0_n_32_622), .A(
      multiplier_0_n_32_621), .B(multiplier_0_n_32_117));
  NAND2_X1_LVT multiplier_0_i_32_147 (.ZN(multiplier_0_n_32_147), .A1(
      multiplier_0_op2_xp[8]), .A2(multiplier_0_op1[11]));
  NAND2_X1_LVT multiplier_0_i_32_131 (.ZN(multiplier_0_n_32_131), .A1(
      multiplier_0_op2_xp[7]), .A2(multiplier_0_op1[12]));
  INV_X1_LVT multiplier_0_i_32_531 (.ZN(multiplier_0_n_32_583), .A(
      multiplier_0_n_32_131));
  NAND2_X1_LVT multiplier_0_i_32_530 (.ZN(multiplier_0_n_32_582), .A1(
      multiplier_0_n_32_147), .A2(multiplier_0_n_32_583));
  NAND2_X1_LVT multiplier_0_i_32_115 (.ZN(multiplier_0_n_32_115), .A1(
      multiplier_0_op2_xp[6]), .A2(multiplier_0_op1[13]));
  INV_X1_LVT multiplier_0_i_32_533 (.ZN(multiplier_0_n_32_585), .A(
      multiplier_0_n_32_115));
  NAND2_X1_LVT multiplier_0_i_32_532 (.ZN(multiplier_0_n_32_584), .A1(
      multiplier_0_n_32_147), .A2(multiplier_0_n_32_585));
  OR2_X1_LVT multiplier_0_i_32_534 (.ZN(multiplier_0_n_32_586), .A1(
      multiplier_0_n_32_115), .A2(multiplier_0_n_32_131));
  NAND3_X1_LVT multiplier_0_i_32_529 (.ZN(multiplier_0_n_32_581), .A1(
      multiplier_0_n_32_582), .A2(multiplier_0_n_32_584), .A3(
      multiplier_0_n_32_586));
  NAND2_X1_LVT multiplier_0_i_32_82 (.ZN(multiplier_0_n_32_82), .A1(
      multiplier_0_op2_xp[4]), .A2(multiplier_0_op1[14]));
  NAND2_X1_LVT multiplier_0_i_32_98 (.ZN(multiplier_0_n_32_98), .A1(
      multiplier_0_op2_xp[5]), .A2(multiplier_0_op1[13]));
  NOR2_X1_LVT multiplier_0_i_32_520 (.ZN(multiplier_0_n_32_568), .A1(
      multiplier_0_n_32_82), .A2(multiplier_0_n_32_98));
  NAND2_X1_LVT multiplier_0_i_32_66 (.ZN(multiplier_0_n_32_66), .A1(
      multiplier_0_op2_xp[3]), .A2(multiplier_0_op1[15]));
  NOR2_X1_LVT multiplier_0_i_32_521 (.ZN(multiplier_0_n_32_569), .A1(
      multiplier_0_n_32_66), .A2(multiplier_0_n_32_98));
  NOR2_X1_LVT multiplier_0_i_32_522 (.ZN(multiplier_0_n_32_570), .A1(
      multiplier_0_n_32_66), .A2(multiplier_0_n_32_82));
  OR3_X1_LVT multiplier_0_i_32_519 (.ZN(multiplier_0_n_32_567), .A1(
      multiplier_0_n_32_568), .A2(multiplier_0_n_32_569), .A3(
      multiplier_0_n_32_570));
  NAND2_X1_LVT multiplier_0_i_32_146 (.ZN(multiplier_0_n_32_146), .A1(
      multiplier_0_op2_xp[8]), .A2(multiplier_0_op1[10]));
  NAND2_X1_LVT multiplier_0_i_32_130 (.ZN(multiplier_0_n_32_130), .A1(
      multiplier_0_op2_xp[7]), .A2(multiplier_0_op1[11]));
  INV_X1_LVT multiplier_0_i_32_512 (.ZN(multiplier_0_n_32_560), .A(
      multiplier_0_n_32_130));
  NAND2_X1_LVT multiplier_0_i_32_511 (.ZN(multiplier_0_n_32_559), .A1(
      multiplier_0_n_32_146), .A2(multiplier_0_n_32_560));
  NAND2_X1_LVT multiplier_0_i_32_114 (.ZN(multiplier_0_n_32_114), .A1(
      multiplier_0_op2_xp[6]), .A2(multiplier_0_op1[12]));
  INV_X1_LVT multiplier_0_i_32_514 (.ZN(multiplier_0_n_32_562), .A(
      multiplier_0_n_32_114));
  NAND2_X1_LVT multiplier_0_i_32_513 (.ZN(multiplier_0_n_32_561), .A1(
      multiplier_0_n_32_146), .A2(multiplier_0_n_32_562));
  OR2_X1_LVT multiplier_0_i_32_515 (.ZN(multiplier_0_n_32_563), .A1(
      multiplier_0_n_32_114), .A2(multiplier_0_n_32_130));
  NAND3_X1_LVT multiplier_0_i_32_510 (.ZN(multiplier_0_n_32_558), .A1(
      multiplier_0_n_32_559), .A2(multiplier_0_n_32_561), .A3(
      multiplier_0_n_32_563));
  NAND2_X1_LVT multiplier_0_i_32_50 (.ZN(multiplier_0_n_32_50), .A1(
      multiplier_0_op2_xp[2]), .A2(multiplier_0_op1_xp[16]));
  NAND2_X1_LVT multiplier_0_i_32_81 (.ZN(multiplier_0_n_32_81), .A1(
      multiplier_0_op2_xp[4]), .A2(multiplier_0_op1[13]));
  NAND2_X1_LVT multiplier_0_i_32_97 (.ZN(multiplier_0_n_32_97), .A1(
      multiplier_0_op2_xp[5]), .A2(multiplier_0_op1[12]));
  NOR2_X1_LVT multiplier_0_i_32_493 (.ZN(multiplier_0_n_32_537), .A1(
      multiplier_0_n_32_81), .A2(multiplier_0_n_32_97));
  NAND2_X1_LVT multiplier_0_i_32_65 (.ZN(multiplier_0_n_32_65), .A1(
      multiplier_0_op2_xp[3]), .A2(multiplier_0_op1[14]));
  NOR2_X1_LVT multiplier_0_i_32_494 (.ZN(multiplier_0_n_32_538), .A1(
      multiplier_0_n_32_65), .A2(multiplier_0_n_32_97));
  NOR2_X1_LVT multiplier_0_i_32_495 (.ZN(multiplier_0_n_32_539), .A1(
      multiplier_0_n_32_65), .A2(multiplier_0_n_32_81));
  OR3_X1_LVT multiplier_0_i_32_492 (.ZN(multiplier_0_n_32_536), .A1(
      multiplier_0_n_32_537), .A2(multiplier_0_n_32_538), .A3(
      multiplier_0_n_32_539));
  NAND2_X1_LVT multiplier_0_i_32_145 (.ZN(multiplier_0_n_32_145), .A1(
      multiplier_0_op2_xp[8]), .A2(multiplier_0_op1[9]));
  NAND2_X1_LVT multiplier_0_i_32_129 (.ZN(multiplier_0_n_32_129), .A1(
      multiplier_0_op2_xp[7]), .A2(multiplier_0_op1[10]));
  INV_X1_LVT multiplier_0_i_32_485 (.ZN(multiplier_0_n_32_529), .A(
      multiplier_0_n_32_129));
  NAND2_X1_LVT multiplier_0_i_32_484 (.ZN(multiplier_0_n_32_528), .A1(
      multiplier_0_n_32_145), .A2(multiplier_0_n_32_529));
  NAND2_X1_LVT multiplier_0_i_32_113 (.ZN(multiplier_0_n_32_113), .A1(
      multiplier_0_op2_xp[6]), .A2(multiplier_0_op1[11]));
  INV_X1_LVT multiplier_0_i_32_487 (.ZN(multiplier_0_n_32_531), .A(
      multiplier_0_n_32_113));
  NAND2_X1_LVT multiplier_0_i_32_486 (.ZN(multiplier_0_n_32_530), .A1(
      multiplier_0_n_32_145), .A2(multiplier_0_n_32_531));
  OR2_X1_LVT multiplier_0_i_32_488 (.ZN(multiplier_0_n_32_532), .A1(
      multiplier_0_n_32_113), .A2(multiplier_0_n_32_129));
  NAND3_X1_LVT multiplier_0_i_32_483 (.ZN(multiplier_0_n_32_527), .A1(
      multiplier_0_n_32_528), .A2(multiplier_0_n_32_530), .A3(
      multiplier_0_n_32_532));
  FA_X1_LVT multiplier_0_i_32_523 (.CO(multiplier_0_n_32_572), .S(
      multiplier_0_n_32_571), .A(multiplier_0_n_32_50), .B(multiplier_0_n_32_536), 
      .CI(multiplier_0_n_32_527));
  FA_X1_LVT multiplier_0_i_32_543 (.CO(multiplier_0_n_32_596), .S(
      multiplier_0_n_32_595), .A(multiplier_0_n_32_567), .B(
      multiplier_0_n_32_558), .CI(multiplier_0_n_32_572));
  XNOR2_X1_LVT multiplier_0_i_32_554 (.ZN(multiplier_0_n_32_609), .A(
      multiplier_0_n_32_100), .B(multiplier_0_n_32_84));
  XNOR2_X1_LVT multiplier_0_i_32_555 (.ZN(multiplier_0_n_32_610), .A(
      multiplier_0_n_32_609), .B(multiplier_0_n_32_589));
  INV_X1_LVT multiplier_0_i_32_556 (.ZN(multiplier_0_n_32_611), .A(
      multiplier_0_n_32_610));
  FA_X1_LVT multiplier_0_i_32_562 (.CO(multiplier_0_n_32_618), .S(
      multiplier_0_n_32_617), .A(multiplier_0_n_32_581), .B(
      multiplier_0_n_32_596), .CI(multiplier_0_n_32_611));
  FA_X1_LVT multiplier_0_i_32_573 (.CO(multiplier_0_n_32_632), .S(
      multiplier_0_n_32_631), .A(multiplier_0_n_32_622), .B(
      multiplier_0_n_32_629), .CI(multiplier_0_n_32_618));
  XNOR2_X1_LVT multiplier_0_i_32_546 (.ZN(multiplier_0_n_32_601), .A(
      multiplier_0_n_32_148), .B(multiplier_0_n_32_132));
  XNOR2_X1_LVT multiplier_0_i_32_547 (.ZN(multiplier_0_n_32_602), .A(
      multiplier_0_n_32_601), .B(multiplier_0_n_32_116));
  XNOR2_X1_LVT multiplier_0_i_32_535 (.ZN(multiplier_0_n_32_587), .A(
      multiplier_0_n_32_99), .B(multiplier_0_n_32_83));
  XNOR2_X1_LVT multiplier_0_i_32_536 (.ZN(multiplier_0_n_32_588), .A(
      multiplier_0_n_32_587), .B(multiplier_0_n_32_67));
  XNOR2_X1_LVT multiplier_0_i_32_527 (.ZN(multiplier_0_n_32_579), .A(
      multiplier_0_n_32_147), .B(multiplier_0_n_32_131));
  XNOR2_X1_LVT multiplier_0_i_32_528 (.ZN(multiplier_0_n_32_580), .A(
      multiplier_0_n_32_579), .B(multiplier_0_n_32_115));
  FA_X1_LVT multiplier_0_i_32_544 (.CO(multiplier_0_n_32_598), .S(
      multiplier_0_n_32_597), .A(multiplier_0_n_32_588), .B(
      multiplier_0_n_32_580), .CI(multiplier_0_n_32_595));
  FA_X1_LVT multiplier_0_i_32_563 (.CO(multiplier_0_n_32_620), .S(
      multiplier_0_n_32_619), .A(multiplier_0_n_32_602), .B(
      multiplier_0_n_32_598), .CI(multiplier_0_n_32_617));
  NAND2_X1_LVT multiplier_0_i_32_33 (.ZN(multiplier_0_n_32_33), .A1(
      multiplier_0_op2_xp[1]), .A2(multiplier_0_op1_xp[16]));
  NAND2_X1_LVT multiplier_0_i_32_49 (.ZN(multiplier_0_n_32_49), .A1(
      multiplier_0_op2_xp[2]), .A2(multiplier_0_op1[15]));
  INV_X1_LVT multiplier_0_i_32_501 (.ZN(multiplier_0_n_32_545), .A(
      multiplier_0_n_32_49));
  NAND2_X1_LVT multiplier_0_i_32_500 (.ZN(multiplier_0_n_32_544), .A1(
      multiplier_0_n_32_33), .A2(multiplier_0_n_32_545));
  NAND2_X1_LVT multiplier_0_i_32_48 (.ZN(multiplier_0_n_32_48), .A1(
      multiplier_0_op2_xp[2]), .A2(multiplier_0_op1[14]));
  NAND2_X1_LVT multiplier_0_i_32_64 (.ZN(multiplier_0_n_32_64), .A1(
      multiplier_0_op2_xp[3]), .A2(multiplier_0_op1[13]));
  NOR2_X1_LVT multiplier_0_i_32_473 (.ZN(multiplier_0_n_32_512), .A1(
      multiplier_0_n_32_48), .A2(multiplier_0_n_32_64));
  NAND2_X1_LVT multiplier_0_i_32_32 (.ZN(multiplier_0_n_32_32), .A1(
      multiplier_0_op2_xp[1]), .A2(multiplier_0_op1[15]));
  NOR2_X1_LVT multiplier_0_i_32_474 (.ZN(multiplier_0_n_32_513), .A1(
      multiplier_0_n_32_32), .A2(multiplier_0_n_32_64));
  NOR2_X1_LVT multiplier_0_i_32_475 (.ZN(multiplier_0_n_32_514), .A1(
      multiplier_0_n_32_32), .A2(multiplier_0_n_32_48));
  OR3_X1_LVT multiplier_0_i_32_472 (.ZN(multiplier_0_n_32_511), .A1(
      multiplier_0_n_32_512), .A2(multiplier_0_n_32_513), .A3(
      multiplier_0_n_32_514));
  NAND2_X1_LVT multiplier_0_i_32_502 (.ZN(multiplier_0_n_32_546), .A1(
      multiplier_0_n_32_511), .A2(multiplier_0_n_32_545));
  NAND2_X1_LVT multiplier_0_i_32_503 (.ZN(multiplier_0_n_32_547), .A1(
      multiplier_0_n_32_511), .A2(multiplier_0_n_32_33));
  NAND3_X1_LVT multiplier_0_i_32_499 (.ZN(multiplier_0_n_32_543), .A1(
      multiplier_0_n_32_544), .A2(multiplier_0_n_32_546), .A3(
      multiplier_0_n_32_547));
  NAND2_X1_LVT multiplier_0_i_32_96 (.ZN(multiplier_0_n_32_96), .A1(
      multiplier_0_op2_xp[5]), .A2(multiplier_0_op1[11]));
  NAND2_X1_LVT multiplier_0_i_32_112 (.ZN(multiplier_0_n_32_112), .A1(
      multiplier_0_op2_xp[6]), .A2(multiplier_0_op1[10]));
  NOR2_X1_LVT multiplier_0_i_32_466 (.ZN(multiplier_0_n_32_505), .A1(
      multiplier_0_n_32_96), .A2(multiplier_0_n_32_112));
  NAND2_X1_LVT multiplier_0_i_32_80 (.ZN(multiplier_0_n_32_80), .A1(
      multiplier_0_op2_xp[4]), .A2(multiplier_0_op1[12]));
  NOR2_X1_LVT multiplier_0_i_32_467 (.ZN(multiplier_0_n_32_506), .A1(
      multiplier_0_n_32_80), .A2(multiplier_0_n_32_112));
  NOR2_X1_LVT multiplier_0_i_32_468 (.ZN(multiplier_0_n_32_507), .A1(
      multiplier_0_n_32_80), .A2(multiplier_0_n_32_96));
  OR3_X1_LVT multiplier_0_i_32_465 (.ZN(multiplier_0_n_32_504), .A1(
      multiplier_0_n_32_505), .A2(multiplier_0_n_32_506), .A3(
      multiplier_0_n_32_507));
  NAND2_X1_LVT multiplier_0_i_32_128 (.ZN(multiplier_0_n_32_128), .A1(
      multiplier_0_op2_xp[7]), .A2(multiplier_0_op1[9]));
  NAND2_X1_LVT multiplier_0_i_32_144 (.ZN(multiplier_0_n_32_144), .A1(
      multiplier_0_op2_xp[8]), .A2(multiplier_0_op1[8]));
  INV_X1_LVT multiplier_0_i_32_461 (.ZN(multiplier_0_n_32_500), .A(
      multiplier_0_n_32_144));
  NAND2_X1_LVT multiplier_0_i_32_460 (.ZN(multiplier_0_n_32_499), .A1(
      multiplier_0_n_32_128), .A2(multiplier_0_n_32_500));
  NAND2_X1_LVT multiplier_0_i_32_16 (.ZN(multiplier_0_n_32_16), .A1(
      multiplier_0_op2_xp[0]), .A2(multiplier_0_op1_xp[16]));
  NOR2_X1_LVT multiplier_0_i_32_451 (.ZN(multiplier_0_n_32_486), .A1(
      multiplier_0_n_32_31), .A2(multiplier_0_n_32_47));
  NOR2_X1_LVT multiplier_0_i_32_452 (.ZN(multiplier_0_n_32_487), .A1(
      multiplier_0_n_32_15), .A2(multiplier_0_n_32_47));
  NOR2_X1_LVT multiplier_0_i_32_453 (.ZN(multiplier_0_n_32_488), .A1(
      multiplier_0_n_32_15), .A2(multiplier_0_n_32_31));
  OR3_X1_LVT multiplier_0_i_32_450 (.ZN(multiplier_0_n_32_485), .A1(
      multiplier_0_n_32_486), .A2(multiplier_0_n_32_487), .A3(
      multiplier_0_n_32_488));
  NOR2_X1_LVT multiplier_0_i_32_444 (.ZN(multiplier_0_n_32_479), .A1(
      multiplier_0_n_32_79), .A2(multiplier_0_n_32_95));
  NOR2_X1_LVT multiplier_0_i_32_445 (.ZN(multiplier_0_n_32_480), .A1(
      multiplier_0_n_32_63), .A2(multiplier_0_n_32_95));
  NOR2_X1_LVT multiplier_0_i_32_446 (.ZN(multiplier_0_n_32_481), .A1(
      multiplier_0_n_32_63), .A2(multiplier_0_n_32_79));
  OR3_X1_LVT multiplier_0_i_32_443 (.ZN(multiplier_0_n_32_478), .A1(
      multiplier_0_n_32_479), .A2(multiplier_0_n_32_480), .A3(
      multiplier_0_n_32_481));
  FA_X1_LVT multiplier_0_i_32_476 (.CO(multiplier_0_n_32_516), .S(
      multiplier_0_n_32_515), .A(multiplier_0_n_32_16), .B(multiplier_0_n_32_485), 
      .CI(multiplier_0_n_32_478));
  FA_X1_LVT multiplier_0_i_32_504 (.CO(multiplier_0_n_32_549), .S(
      multiplier_0_n_32_548), .A(multiplier_0_n_32_504), .B(
      multiplier_0_n_32_499), .CI(multiplier_0_n_32_516));
  XNOR2_X1_LVT multiplier_0_i_32_516 (.ZN(multiplier_0_n_32_564), .A(
      multiplier_0_n_32_98), .B(multiplier_0_n_32_82));
  XNOR2_X1_LVT multiplier_0_i_32_517 (.ZN(multiplier_0_n_32_565), .A(
      multiplier_0_n_32_564), .B(multiplier_0_n_32_66));
  INV_X1_LVT multiplier_0_i_32_518 (.ZN(multiplier_0_n_32_566), .A(
      multiplier_0_n_32_565));
  FA_X1_LVT multiplier_0_i_32_524 (.CO(multiplier_0_n_32_574), .S(
      multiplier_0_n_32_573), .A(multiplier_0_n_32_543), .B(
      multiplier_0_n_32_549), .CI(multiplier_0_n_32_566));
  XNOR2_X1_LVT multiplier_0_i_32_508 (.ZN(multiplier_0_n_32_556), .A(
      multiplier_0_n_32_146), .B(multiplier_0_n_32_130));
  XNOR2_X1_LVT multiplier_0_i_32_509 (.ZN(multiplier_0_n_32_557), .A(
      multiplier_0_n_32_556), .B(multiplier_0_n_32_114));
  XNOR2_X1_LVT multiplier_0_i_32_496 (.ZN(multiplier_0_n_32_540), .A(
      multiplier_0_n_32_49), .B(multiplier_0_n_32_33));
  XNOR2_X1_LVT multiplier_0_i_32_497 (.ZN(multiplier_0_n_32_541), .A(
      multiplier_0_n_32_540), .B(multiplier_0_n_32_511));
  INV_X1_LVT multiplier_0_i_32_498 (.ZN(multiplier_0_n_32_542), .A(
      multiplier_0_n_32_541));
  XNOR2_X1_LVT multiplier_0_i_32_489 (.ZN(multiplier_0_n_32_533), .A(
      multiplier_0_n_32_97), .B(multiplier_0_n_32_81));
  XNOR2_X1_LVT multiplier_0_i_32_490 (.ZN(multiplier_0_n_32_534), .A(
      multiplier_0_n_32_533), .B(multiplier_0_n_32_65));
  INV_X1_LVT multiplier_0_i_32_491 (.ZN(multiplier_0_n_32_535), .A(
      multiplier_0_n_32_534));
  XNOR2_X1_LVT multiplier_0_i_32_481 (.ZN(multiplier_0_n_32_525), .A(
      multiplier_0_n_32_145), .B(multiplier_0_n_32_129));
  XNOR2_X1_LVT multiplier_0_i_32_482 (.ZN(multiplier_0_n_32_526), .A(
      multiplier_0_n_32_525), .B(multiplier_0_n_32_113));
  FA_X1_LVT multiplier_0_i_32_505 (.CO(multiplier_0_n_32_551), .S(
      multiplier_0_n_32_550), .A(multiplier_0_n_32_542), .B(
      multiplier_0_n_32_535), .CI(multiplier_0_n_32_526));
  FA_X1_LVT multiplier_0_i_32_525 (.CO(multiplier_0_n_32_576), .S(
      multiplier_0_n_32_575), .A(multiplier_0_n_32_557), .B(
      multiplier_0_n_32_571), .CI(multiplier_0_n_32_551));
  FA_X1_LVT multiplier_0_i_32_545 (.CO(multiplier_0_n_32_600), .S(
      multiplier_0_n_32_599), .A(multiplier_0_n_32_574), .B(
      multiplier_0_n_32_576), .CI(multiplier_0_n_32_597));
  INV_X1_LVT multiplier_0_i_32_436 (.ZN(multiplier_0_n_32_471), .A(
      multiplier_0_n_32_127));
  NAND2_X1_LVT multiplier_0_i_32_435 (.ZN(multiplier_0_n_32_470), .A1(
      multiplier_0_n_32_143), .A2(multiplier_0_n_32_471));
  INV_X1_LVT multiplier_0_i_32_438 (.ZN(multiplier_0_n_32_473), .A(
      multiplier_0_n_32_111));
  NAND2_X1_LVT multiplier_0_i_32_437 (.ZN(multiplier_0_n_32_472), .A1(
      multiplier_0_n_32_143), .A2(multiplier_0_n_32_473));
  OR2_X1_LVT multiplier_0_i_32_439 (.ZN(multiplier_0_n_32_474), .A1(
      multiplier_0_n_32_111), .A2(multiplier_0_n_32_127));
  NAND3_X1_LVT multiplier_0_i_32_434 (.ZN(multiplier_0_n_32_469), .A1(
      multiplier_0_n_32_470), .A2(multiplier_0_n_32_472), .A3(
      multiplier_0_n_32_474));
  XNOR2_X1_LVT multiplier_0_i_32_469 (.ZN(multiplier_0_n_32_508), .A(
      multiplier_0_n_32_64), .B(multiplier_0_n_32_48));
  XNOR2_X1_LVT multiplier_0_i_32_470 (.ZN(multiplier_0_n_32_509), .A(
      multiplier_0_n_32_508), .B(multiplier_0_n_32_32));
  INV_X1_LVT multiplier_0_i_32_471 (.ZN(multiplier_0_n_32_510), .A(
      multiplier_0_n_32_509));
  FA_X1_LVT multiplier_0_i_32_477 (.CO(multiplier_0_n_32_518), .S(
      multiplier_0_n_32_517), .A(multiplier_0_n_32_469), .B(
      multiplier_0_n_32_490), .CI(multiplier_0_n_32_510));
  XNOR2_X1_LVT multiplier_0_i_32_462 (.ZN(multiplier_0_n_32_501), .A(
      multiplier_0_n_32_112), .B(multiplier_0_n_32_96));
  XNOR2_X1_LVT multiplier_0_i_32_463 (.ZN(multiplier_0_n_32_502), .A(
      multiplier_0_n_32_501), .B(multiplier_0_n_32_80));
  INV_X1_LVT multiplier_0_i_32_464 (.ZN(multiplier_0_n_32_503), .A(
      multiplier_0_n_32_502));
  XNOR2_X1_LVT multiplier_0_i_32_458 (.ZN(multiplier_0_n_32_497), .A(
      multiplier_0_n_32_144), .B(multiplier_0_n_32_128));
  INV_X1_LVT multiplier_0_i_32_459 (.ZN(multiplier_0_n_32_498), .A(
      multiplier_0_n_32_497));
  FA_X1_LVT multiplier_0_i_32_478 (.CO(multiplier_0_n_32_520), .S(
      multiplier_0_n_32_519), .A(multiplier_0_n_32_503), .B(
      multiplier_0_n_32_498), .CI(multiplier_0_n_32_515));
  FA_X1_LVT multiplier_0_i_32_506 (.CO(multiplier_0_n_32_553), .S(
      multiplier_0_n_32_552), .A(multiplier_0_n_32_548), .B(
      multiplier_0_n_32_518), .CI(multiplier_0_n_32_520));
  FA_X1_LVT multiplier_0_i_32_526 (.CO(multiplier_0_n_32_578), .S(
      multiplier_0_n_32_577), .A(multiplier_0_n_32_573), .B(
      multiplier_0_n_32_553), .CI(multiplier_0_n_32_575));
  FA_X1_LVT multiplier_0_i_32_479 (.CO(multiplier_0_n_32_522), .S(
      multiplier_0_n_32_521), .A(multiplier_0_n_32_492), .B(
      multiplier_0_n_32_517), .CI(multiplier_0_n_32_494));
  FA_X1_LVT multiplier_0_i_32_507 (.CO(multiplier_0_n_32_555), .S(
      multiplier_0_n_32_554), .A(multiplier_0_n_32_522), .B(
      multiplier_0_n_32_550), .CI(multiplier_0_n_32_552));
  HA_X1_LVT multiplier_0_i_32_480 (.CO(multiplier_0_n_32_524), .S(
      multiplier_0_n_32_523), .A(multiplier_0_n_32_519), .B(
      multiplier_0_n_32_521));
  FA_X1_LVT multiplier_0_i_32_610 (.CO(multiplier_0_n_32_667), .S(
      multiplier_0_n_58), .A(multiplier_0_n_32_496), .B(multiplier_0_n_32_523), 
      .CI(multiplier_0_n_32_666));
  FA_X1_LVT multiplier_0_i_32_611 (.CO(multiplier_0_n_32_668), .S(
      multiplier_0_n_59), .A(multiplier_0_n_32_524), .B(multiplier_0_n_32_554), 
      .CI(multiplier_0_n_32_667));
  FA_X1_LVT multiplier_0_i_32_612 (.CO(multiplier_0_n_32_669), .S(
      multiplier_0_n_60), .A(multiplier_0_n_32_555), .B(multiplier_0_n_32_577), 
      .CI(multiplier_0_n_32_668));
  FA_X1_LVT multiplier_0_i_32_613 (.CO(multiplier_0_n_32_670), .S(
      multiplier_0_n_61), .A(multiplier_0_n_32_599), .B(multiplier_0_n_32_578), 
      .CI(multiplier_0_n_32_669));
  FA_X1_LVT multiplier_0_i_32_614 (.CO(multiplier_0_n_32_671), .S(
      multiplier_0_n_62), .A(multiplier_0_n_32_600), .B(multiplier_0_n_32_619), 
      .CI(multiplier_0_n_32_670));
  FA_X1_LVT multiplier_0_i_32_615 (.CO(multiplier_0_n_32_672), .S(
      multiplier_0_n_63), .A(multiplier_0_n_32_620), .B(multiplier_0_n_32_631), 
      .CI(multiplier_0_n_32_671));
  FA_X1_LVT multiplier_0_i_32_616 (.CO(multiplier_0_n_32_673), .S(
      multiplier_0_n_64), .A(multiplier_0_n_32_632), .B(multiplier_0_n_32_641), 
      .CI(multiplier_0_n_32_672));
  XNOR2_X1_LVT multiplier_0_i_32_618 (.ZN(multiplier_0_n_65), .A(
      multiplier_0_n_32_674), .B(multiplier_0_n_32_673));
  AND2_X1_LVT multiplier_0_i_33_0 (.ZN(multiplier_0_n_66), .A1(
      multiplier_0_sign_sel), .A2(multiplier_0_n_65));
  NAND2_X1_LVT multiplier_0_i_34_49 (.ZN(multiplier_0_n_34_25), .A1(
      multiplier_0_n_34_8), .A2(multiplier_0_n_66));
  INV_X1_LVT multiplier_0_i_34_47 (.ZN(multiplier_0_n_34_24), .A(
      multiplier_0_n_65));
  OAI21_X1_LVT multiplier_0_i_34_57 (.ZN(multiplier_0_product_xp[31]), .A(
      multiplier_0_n_34_25), .B1(multiplier_0_n_34_8), .B2(multiplier_0_n_34_24));
  NOR3_X1_LVT multiplier_0_i_3_9 (.ZN(multiplier_0_n_7), .A1(multiplier_0_n_3_2), 
      .A2(multiplier_0_n_3_1), .A3(per_addr[0]));
  AND2_X1_LVT multiplier_0_i_7_6 (.ZN(multiplier_0_reshi_wr), .A1(
      multiplier_0_reg_write), .A2(multiplier_0_n_7));
  NOR2_X1_LVT multiplier_0_i_41_0 (.ZN(multiplier_0_n_41_0), .A1(
      multiplier_0_result_clr), .A2(multiplier_0_reshi_wr));
  AOI22_X1_LVT multiplier_0_i_41_31 (.ZN(multiplier_0_n_41_16), .A1(
      multiplier_0_n_41_0), .A2(multiplier_0_reshi_nxt[15]), .B1(
      multiplier_0_reshi_wr), .B2(multiplier_0_per_din_msk[15]));
  INV_X1_LVT multiplier_0_i_41_32 (.ZN(multiplier_0_n_86), .A(
      multiplier_0_n_41_16));
  INV_X1_LVT multiplier_0_i_42_1 (.ZN(multiplier_0_n_42_1), .A(multiplier_0_n_69));
  INV_X1_LVT multiplier_0_i_42_0 (.ZN(multiplier_0_n_42_0), .A(
      multiplier_0_reshi_wr));
  NAND2_X1_LVT multiplier_0_i_42_2 (.ZN(multiplier_0_n_87), .A1(
      multiplier_0_n_42_1), .A2(multiplier_0_n_42_0));
  CLKGATETST_X1_LVT multiplier_0_clk_gate_reshi_reg (.GCK(multiplier_0_n_70), 
      .CK(mclk), .E(multiplier_0_n_87), .SE(1'b0));
  DFFR_X1_LVT \multiplier_0_reshi_reg[15] (.Q(multiplier_0_reshi[15]), .QN(), 
      .CK(multiplier_0_n_70), .D(multiplier_0_n_86), .RN(multiplier_0_n_38));
  INV_X1_LVT multiplier_0_i_34_45 (.ZN(multiplier_0_n_34_23), .A(
      multiplier_0_n_64));
  OAI21_X1_LVT multiplier_0_i_34_56 (.ZN(multiplier_0_product_xp[30]), .A(
      multiplier_0_n_34_25), .B1(multiplier_0_n_34_8), .B2(multiplier_0_n_34_23));
  AOI22_X1_LVT multiplier_0_i_41_29 (.ZN(multiplier_0_n_41_15), .A1(
      multiplier_0_n_41_0), .A2(multiplier_0_reshi_nxt[14]), .B1(
      multiplier_0_reshi_wr), .B2(multiplier_0_per_din_msk[14]));
  INV_X1_LVT multiplier_0_i_41_30 (.ZN(multiplier_0_n_85), .A(
      multiplier_0_n_41_15));
  DFFR_X1_LVT \multiplier_0_reshi_reg[14] (.Q(multiplier_0_reshi[14]), .QN(), 
      .CK(multiplier_0_n_70), .D(multiplier_0_n_85), .RN(multiplier_0_n_38));
  INV_X1_LVT multiplier_0_i_34_43 (.ZN(multiplier_0_n_34_22), .A(
      multiplier_0_n_63));
  OAI21_X1_LVT multiplier_0_i_34_55 (.ZN(multiplier_0_product_xp[29]), .A(
      multiplier_0_n_34_25), .B1(multiplier_0_n_34_8), .B2(multiplier_0_n_34_22));
  AOI22_X1_LVT multiplier_0_i_41_27 (.ZN(multiplier_0_n_41_14), .A1(
      multiplier_0_n_41_0), .A2(multiplier_0_reshi_nxt[13]), .B1(
      multiplier_0_reshi_wr), .B2(multiplier_0_per_din_msk[13]));
  INV_X1_LVT multiplier_0_i_41_28 (.ZN(multiplier_0_n_84), .A(
      multiplier_0_n_41_14));
  DFFR_X1_LVT \multiplier_0_reshi_reg[13] (.Q(multiplier_0_reshi[13]), .QN(), 
      .CK(multiplier_0_n_70), .D(multiplier_0_n_84), .RN(multiplier_0_n_38));
  INV_X1_LVT multiplier_0_i_34_41 (.ZN(multiplier_0_n_34_21), .A(
      multiplier_0_n_62));
  OAI21_X1_LVT multiplier_0_i_34_54 (.ZN(multiplier_0_product_xp[28]), .A(
      multiplier_0_n_34_25), .B1(multiplier_0_n_34_8), .B2(multiplier_0_n_34_21));
  AOI22_X1_LVT multiplier_0_i_41_25 (.ZN(multiplier_0_n_41_13), .A1(
      multiplier_0_n_41_0), .A2(multiplier_0_reshi_nxt[12]), .B1(
      multiplier_0_reshi_wr), .B2(multiplier_0_per_din_msk[12]));
  INV_X1_LVT multiplier_0_i_41_26 (.ZN(multiplier_0_n_83), .A(
      multiplier_0_n_41_13));
  DFFR_X1_LVT \multiplier_0_reshi_reg[12] (.Q(multiplier_0_reshi[12]), .QN(), 
      .CK(multiplier_0_n_70), .D(multiplier_0_n_83), .RN(multiplier_0_n_38));
  INV_X1_LVT multiplier_0_i_34_39 (.ZN(multiplier_0_n_34_20), .A(
      multiplier_0_n_61));
  OAI21_X1_LVT multiplier_0_i_34_53 (.ZN(multiplier_0_product_xp[27]), .A(
      multiplier_0_n_34_25), .B1(multiplier_0_n_34_8), .B2(multiplier_0_n_34_20));
  AOI22_X1_LVT multiplier_0_i_41_23 (.ZN(multiplier_0_n_41_12), .A1(
      multiplier_0_n_41_0), .A2(multiplier_0_reshi_nxt[11]), .B1(
      multiplier_0_reshi_wr), .B2(multiplier_0_per_din_msk[11]));
  INV_X1_LVT multiplier_0_i_41_24 (.ZN(multiplier_0_n_82), .A(
      multiplier_0_n_41_12));
  DFFR_X1_LVT \multiplier_0_reshi_reg[11] (.Q(multiplier_0_reshi[11]), .QN(), 
      .CK(multiplier_0_n_70), .D(multiplier_0_n_82), .RN(multiplier_0_n_38));
  INV_X1_LVT multiplier_0_i_34_37 (.ZN(multiplier_0_n_34_19), .A(
      multiplier_0_n_60));
  OAI21_X1_LVT multiplier_0_i_34_52 (.ZN(multiplier_0_product_xp[26]), .A(
      multiplier_0_n_34_25), .B1(multiplier_0_n_34_8), .B2(multiplier_0_n_34_19));
  AOI22_X1_LVT multiplier_0_i_41_21 (.ZN(multiplier_0_n_41_11), .A1(
      multiplier_0_n_41_0), .A2(multiplier_0_reshi_nxt[10]), .B1(
      multiplier_0_reshi_wr), .B2(multiplier_0_per_din_msk[10]));
  INV_X1_LVT multiplier_0_i_41_22 (.ZN(multiplier_0_n_81), .A(
      multiplier_0_n_41_11));
  DFFR_X1_LVT \multiplier_0_reshi_reg[10] (.Q(multiplier_0_reshi[10]), .QN(), 
      .CK(multiplier_0_n_70), .D(multiplier_0_n_81), .RN(multiplier_0_n_38));
  INV_X1_LVT multiplier_0_i_34_35 (.ZN(multiplier_0_n_34_18), .A(
      multiplier_0_n_59));
  OAI21_X1_LVT multiplier_0_i_34_51 (.ZN(multiplier_0_product_xp[25]), .A(
      multiplier_0_n_34_25), .B1(multiplier_0_n_34_8), .B2(multiplier_0_n_34_18));
  AOI22_X1_LVT multiplier_0_i_41_19 (.ZN(multiplier_0_n_41_10), .A1(
      multiplier_0_n_41_0), .A2(multiplier_0_reshi_nxt[9]), .B1(
      multiplier_0_reshi_wr), .B2(multiplier_0_per_din_msk[9]));
  INV_X1_LVT multiplier_0_i_41_20 (.ZN(multiplier_0_n_80), .A(
      multiplier_0_n_41_10));
  DFFR_X1_LVT \multiplier_0_reshi_reg[9] (.Q(multiplier_0_reshi[9]), .QN(), .CK(
      multiplier_0_n_70), .D(multiplier_0_n_80), .RN(multiplier_0_n_38));
  INV_X1_LVT multiplier_0_i_34_33 (.ZN(multiplier_0_n_34_17), .A(
      multiplier_0_n_58));
  OAI21_X1_LVT multiplier_0_i_34_50 (.ZN(multiplier_0_product_xp[24]), .A(
      multiplier_0_n_34_25), .B1(multiplier_0_n_34_8), .B2(multiplier_0_n_34_17));
  AOI22_X1_LVT multiplier_0_i_41_17 (.ZN(multiplier_0_n_41_9), .A1(
      multiplier_0_n_41_0), .A2(multiplier_0_reshi_nxt[8]), .B1(
      multiplier_0_reshi_wr), .B2(multiplier_0_per_din_msk[8]));
  INV_X1_LVT multiplier_0_i_41_18 (.ZN(multiplier_0_n_79), .A(
      multiplier_0_n_41_9));
  DFFR_X1_LVT \multiplier_0_reshi_reg[8] (.Q(multiplier_0_reshi[8]), .QN(), .CK(
      multiplier_0_n_70), .D(multiplier_0_n_79), .RN(multiplier_0_n_38));
  OAI22_X1_LVT multiplier_0_i_34_48 (.ZN(multiplier_0_product_xp[23]), .A1(
      multiplier_0_n_34_8), .A2(multiplier_0_n_34_16), .B1(multiplier_0_n_34_24), 
      .B2(multiplier_0_cycle[0]));
  AOI22_X1_LVT multiplier_0_i_41_15 (.ZN(multiplier_0_n_41_8), .A1(
      multiplier_0_n_41_0), .A2(multiplier_0_reshi_nxt[7]), .B1(
      multiplier_0_reshi_wr), .B2(per_din[7]));
  INV_X1_LVT multiplier_0_i_41_16 (.ZN(multiplier_0_n_78), .A(
      multiplier_0_n_41_8));
  DFFR_X1_LVT \multiplier_0_reshi_reg[7] (.Q(multiplier_0_reshi[7]), .QN(), .CK(
      multiplier_0_n_70), .D(multiplier_0_n_78), .RN(multiplier_0_n_38));
  OAI22_X1_LVT multiplier_0_i_34_46 (.ZN(multiplier_0_product_xp[22]), .A1(
      multiplier_0_n_34_8), .A2(multiplier_0_n_34_15), .B1(multiplier_0_n_34_23), 
      .B2(multiplier_0_cycle[0]));
  AOI22_X1_LVT multiplier_0_i_41_13 (.ZN(multiplier_0_n_41_7), .A1(
      multiplier_0_n_41_0), .A2(multiplier_0_reshi_nxt[6]), .B1(
      multiplier_0_reshi_wr), .B2(per_din[6]));
  INV_X1_LVT multiplier_0_i_41_14 (.ZN(multiplier_0_n_77), .A(
      multiplier_0_n_41_7));
  DFFR_X1_LVT \multiplier_0_reshi_reg[6] (.Q(multiplier_0_reshi[6]), .QN(), .CK(
      multiplier_0_n_70), .D(multiplier_0_n_77), .RN(multiplier_0_n_38));
  OAI22_X1_LVT multiplier_0_i_34_44 (.ZN(multiplier_0_product_xp[21]), .A1(
      multiplier_0_n_34_8), .A2(multiplier_0_n_34_14), .B1(multiplier_0_n_34_22), 
      .B2(multiplier_0_cycle[0]));
  AOI22_X1_LVT multiplier_0_i_41_11 (.ZN(multiplier_0_n_41_6), .A1(
      multiplier_0_n_41_0), .A2(multiplier_0_reshi_nxt[5]), .B1(
      multiplier_0_reshi_wr), .B2(per_din[5]));
  INV_X1_LVT multiplier_0_i_41_12 (.ZN(multiplier_0_n_76), .A(
      multiplier_0_n_41_6));
  DFFR_X1_LVT \multiplier_0_reshi_reg[5] (.Q(multiplier_0_reshi[5]), .QN(), .CK(
      multiplier_0_n_70), .D(multiplier_0_n_76), .RN(multiplier_0_n_38));
  OAI22_X1_LVT multiplier_0_i_34_42 (.ZN(multiplier_0_product_xp[20]), .A1(
      multiplier_0_n_34_8), .A2(multiplier_0_n_34_13), .B1(multiplier_0_n_34_21), 
      .B2(multiplier_0_cycle[0]));
  AOI22_X1_LVT multiplier_0_i_41_9 (.ZN(multiplier_0_n_41_5), .A1(
      multiplier_0_n_41_0), .A2(multiplier_0_reshi_nxt[4]), .B1(
      multiplier_0_reshi_wr), .B2(per_din[4]));
  INV_X1_LVT multiplier_0_i_41_10 (.ZN(multiplier_0_n_75), .A(
      multiplier_0_n_41_5));
  DFFR_X1_LVT \multiplier_0_reshi_reg[4] (.Q(multiplier_0_reshi[4]), .QN(), .CK(
      multiplier_0_n_70), .D(multiplier_0_n_75), .RN(multiplier_0_n_38));
  OAI22_X1_LVT multiplier_0_i_34_40 (.ZN(multiplier_0_product_xp[19]), .A1(
      multiplier_0_n_34_8), .A2(multiplier_0_n_34_12), .B1(multiplier_0_n_34_20), 
      .B2(multiplier_0_cycle[0]));
  AOI22_X1_LVT multiplier_0_i_41_7 (.ZN(multiplier_0_n_41_4), .A1(
      multiplier_0_n_41_0), .A2(multiplier_0_reshi_nxt[3]), .B1(
      multiplier_0_reshi_wr), .B2(per_din[3]));
  INV_X1_LVT multiplier_0_i_41_8 (.ZN(multiplier_0_n_74), .A(multiplier_0_n_41_4));
  DFFR_X1_LVT \multiplier_0_reshi_reg[3] (.Q(multiplier_0_reshi[3]), .QN(), .CK(
      multiplier_0_n_70), .D(multiplier_0_n_74), .RN(multiplier_0_n_38));
  OAI22_X1_LVT multiplier_0_i_34_38 (.ZN(multiplier_0_product_xp[18]), .A1(
      multiplier_0_n_34_8), .A2(multiplier_0_n_34_11), .B1(multiplier_0_n_34_19), 
      .B2(multiplier_0_cycle[0]));
  AOI22_X1_LVT multiplier_0_i_41_5 (.ZN(multiplier_0_n_41_3), .A1(
      multiplier_0_n_41_0), .A2(multiplier_0_reshi_nxt[2]), .B1(
      multiplier_0_reshi_wr), .B2(per_din[2]));
  INV_X1_LVT multiplier_0_i_41_6 (.ZN(multiplier_0_n_73), .A(multiplier_0_n_41_3));
  DFFR_X1_LVT \multiplier_0_reshi_reg[2] (.Q(multiplier_0_reshi[2]), .QN(), .CK(
      multiplier_0_n_70), .D(multiplier_0_n_73), .RN(multiplier_0_n_38));
  OAI22_X1_LVT multiplier_0_i_34_36 (.ZN(multiplier_0_product_xp[17]), .A1(
      multiplier_0_n_34_8), .A2(multiplier_0_n_34_10), .B1(multiplier_0_n_34_18), 
      .B2(multiplier_0_cycle[0]));
  AOI22_X1_LVT multiplier_0_i_41_3 (.ZN(multiplier_0_n_41_2), .A1(
      multiplier_0_n_41_0), .A2(multiplier_0_reshi_nxt[1]), .B1(
      multiplier_0_reshi_wr), .B2(per_din[1]));
  INV_X1_LVT multiplier_0_i_41_4 (.ZN(multiplier_0_n_72), .A(multiplier_0_n_41_2));
  DFFR_X1_LVT \multiplier_0_reshi_reg[1] (.Q(multiplier_0_reshi[1]), .QN(), .CK(
      multiplier_0_n_70), .D(multiplier_0_n_72), .RN(multiplier_0_n_38));
  OAI22_X1_LVT multiplier_0_i_34_34 (.ZN(multiplier_0_product_xp[16]), .A1(
      multiplier_0_n_34_8), .A2(multiplier_0_n_34_9), .B1(multiplier_0_n_34_17), 
      .B2(multiplier_0_cycle[0]));
  AOI22_X1_LVT multiplier_0_i_41_1 (.ZN(multiplier_0_n_41_1), .A1(
      multiplier_0_n_41_0), .A2(multiplier_0_reshi_nxt[0]), .B1(per_din[0]), .B2(
      multiplier_0_reshi_wr));
  INV_X1_LVT multiplier_0_i_41_2 (.ZN(multiplier_0_n_71), .A(multiplier_0_n_41_1));
  DFFR_X1_LVT \multiplier_0_reshi_reg[0] (.Q(multiplier_0_reshi[0]), .QN(), .CK(
      multiplier_0_n_70), .D(multiplier_0_n_71), .RN(multiplier_0_n_38));
  FA_X1_LVT multiplier_0_i_48_16 (.CO(multiplier_0_n_48_16), .S(
      multiplier_0_reshi_nxt[0]), .A(multiplier_0_product_xp[16]), .B(
      multiplier_0_reshi[0]), .CI(multiplier_0_n_48_15));
  FA_X1_LVT multiplier_0_i_48_17 (.CO(multiplier_0_n_48_17), .S(
      multiplier_0_reshi_nxt[1]), .A(multiplier_0_product_xp[17]), .B(
      multiplier_0_reshi[1]), .CI(multiplier_0_n_48_16));
  FA_X1_LVT multiplier_0_i_48_18 (.CO(multiplier_0_n_48_18), .S(
      multiplier_0_reshi_nxt[2]), .A(multiplier_0_product_xp[18]), .B(
      multiplier_0_reshi[2]), .CI(multiplier_0_n_48_17));
  FA_X1_LVT multiplier_0_i_48_19 (.CO(multiplier_0_n_48_19), .S(
      multiplier_0_reshi_nxt[3]), .A(multiplier_0_product_xp[19]), .B(
      multiplier_0_reshi[3]), .CI(multiplier_0_n_48_18));
  FA_X1_LVT multiplier_0_i_48_20 (.CO(multiplier_0_n_48_20), .S(
      multiplier_0_reshi_nxt[4]), .A(multiplier_0_product_xp[20]), .B(
      multiplier_0_reshi[4]), .CI(multiplier_0_n_48_19));
  FA_X1_LVT multiplier_0_i_48_21 (.CO(multiplier_0_n_48_21), .S(
      multiplier_0_reshi_nxt[5]), .A(multiplier_0_product_xp[21]), .B(
      multiplier_0_reshi[5]), .CI(multiplier_0_n_48_20));
  FA_X1_LVT multiplier_0_i_48_22 (.CO(multiplier_0_n_48_22), .S(
      multiplier_0_reshi_nxt[6]), .A(multiplier_0_product_xp[22]), .B(
      multiplier_0_reshi[6]), .CI(multiplier_0_n_48_21));
  FA_X1_LVT multiplier_0_i_48_23 (.CO(multiplier_0_n_48_23), .S(
      multiplier_0_reshi_nxt[7]), .A(multiplier_0_product_xp[23]), .B(
      multiplier_0_reshi[7]), .CI(multiplier_0_n_48_22));
  FA_X1_LVT multiplier_0_i_48_24 (.CO(multiplier_0_n_48_24), .S(
      multiplier_0_reshi_nxt[8]), .A(multiplier_0_product_xp[24]), .B(
      multiplier_0_reshi[8]), .CI(multiplier_0_n_48_23));
  FA_X1_LVT multiplier_0_i_48_25 (.CO(multiplier_0_n_48_25), .S(
      multiplier_0_reshi_nxt[9]), .A(multiplier_0_product_xp[25]), .B(
      multiplier_0_reshi[9]), .CI(multiplier_0_n_48_24));
  FA_X1_LVT multiplier_0_i_48_26 (.CO(multiplier_0_n_48_26), .S(
      multiplier_0_reshi_nxt[10]), .A(multiplier_0_product_xp[26]), .B(
      multiplier_0_reshi[10]), .CI(multiplier_0_n_48_25));
  FA_X1_LVT multiplier_0_i_48_27 (.CO(multiplier_0_n_48_27), .S(
      multiplier_0_reshi_nxt[11]), .A(multiplier_0_product_xp[27]), .B(
      multiplier_0_reshi[11]), .CI(multiplier_0_n_48_26));
  FA_X1_LVT multiplier_0_i_48_28 (.CO(multiplier_0_n_48_28), .S(
      multiplier_0_reshi_nxt[12]), .A(multiplier_0_product_xp[28]), .B(
      multiplier_0_reshi[12]), .CI(multiplier_0_n_48_27));
  FA_X1_LVT multiplier_0_i_48_29 (.CO(multiplier_0_n_48_29), .S(
      multiplier_0_reshi_nxt[13]), .A(multiplier_0_product_xp[29]), .B(
      multiplier_0_reshi[13]), .CI(multiplier_0_n_48_28));
  FA_X1_LVT multiplier_0_i_48_30 (.CO(multiplier_0_n_48_30), .S(
      multiplier_0_reshi_nxt[14]), .A(multiplier_0_product_xp[30]), .B(
      multiplier_0_reshi[14]), .CI(multiplier_0_n_48_29));
  FA_X1_LVT multiplier_0_i_48_31 (.CO(multiplier_0_n_138), .S(
      multiplier_0_reshi_nxt[15]), .A(multiplier_0_product_xp[31]), .B(
      multiplier_0_reshi[15]), .CI(multiplier_0_n_48_30));
  NAND2_X1_LVT multiplier_0_i_50_0 (.ZN(multiplier_0_n_50_0), .A1(
      multiplier_0_reshi_nxt[15]), .A2(multiplier_0_sign_sel));
  INV_X1_LVT multiplier_0_i_50_3 (.ZN(multiplier_0_sumext_s_nxt[1]), .A(
      multiplier_0_n_50_0));
  AND2_X1_LVT multiplier_0_i_52_2 (.ZN(multiplier_0_n_142), .A1(
      multiplier_0_n_52_0), .A2(multiplier_0_sumext_s_nxt[1]));
  INV_X1_LVT multiplier_0_i_53_1 (.ZN(multiplier_0_n_53_1), .A(
      multiplier_0_result_wr));
  INV_X1_LVT multiplier_0_i_53_0 (.ZN(multiplier_0_n_53_0), .A(
      multiplier_0_op2_wr));
  NAND2_X1_LVT multiplier_0_i_53_2 (.ZN(multiplier_0_n_143), .A1(
      multiplier_0_n_53_1), .A2(multiplier_0_n_53_0));
  CLKGATETST_X1_LVT multiplier_0_clk_gate_sumext_s_reg (.GCK(multiplier_0_n_140), 
      .CK(mclk), .E(multiplier_0_n_143), .SE(1'b0));
  DFFR_X1_LVT \multiplier_0_sumext_s_reg[1] (.Q(multiplier_0_sumext_s[1]), .QN(), 
      .CK(multiplier_0_n_140), .D(multiplier_0_n_142), .RN(multiplier_0_n_38));
  AOI22_X1_LVT multiplier_0_i_57_1 (.ZN(multiplier_0_n_57_1), .A1(
      multiplier_0_n_57_0), .A2(multiplier_0_sumext_s[1]), .B1(
      multiplier_0_sumext_s_nxt[1]), .B2(multiplier_0_cycle[1]));
  INV_X1_LVT multiplier_0_i_57_2 (.ZN(multiplier_0_n_148), .A(
      multiplier_0_n_57_1));
  NOR3_X1_LVT multiplier_0_i_3_10 (.ZN(multiplier_0_n_8), .A1(multiplier_0_n_3_0), 
      .A2(multiplier_0_n_3_1), .A3(multiplier_0_n_3_2));
  AND2_X1_LVT multiplier_0_i_4_7 (.ZN(multiplier_0_reg_rd15), .A1(
      multiplier_0_reg_read), .A2(multiplier_0_n_8));
  AND2_X1_LVT multiplier_0_i_58_0 (.ZN(multiplier_0_n_149), .A1(
      multiplier_0_n_148), .A2(multiplier_0_reg_rd15));
  AND2_X1_LVT multiplier_0_i_4_4 (.ZN(multiplier_0_n_12), .A1(
      multiplier_0_reg_read), .A2(multiplier_0_n_5));
  AND2_X1_LVT multiplier_0_i_20_0 (.ZN(multiplier_0_n_37), .A1(
      multiplier_0_op2_reg[15]), .A2(multiplier_0_n_12));
  NOR4_X1_LVT multiplier_0_i_60_96 (.ZN(multiplier_0_n_60_81), .A1(
      multiplier_0_n_60_79), .A2(multiplier_0_n_60_80), .A3(multiplier_0_n_149), 
      .A4(multiplier_0_n_37));
  AOI22_X1_LVT multiplier_0_i_60_97 (.ZN(multiplier_0_n_60_82), .A1(
      multiplier_0_n_60_0), .A2(multiplier_0_reshi[15]), .B1(
      multiplier_0_cycle[1]), .B2(multiplier_0_reshi_nxt[15]));
  AND2_X1_LVT multiplier_0_i_4_6 (.ZN(multiplier_0_n_14), .A1(
      multiplier_0_reg_read), .A2(multiplier_0_n_7));
  INV_X1_LVT multiplier_0_i_60_7 (.ZN(multiplier_0_n_60_7), .A(multiplier_0_n_14));
  OAI21_X1_LVT multiplier_0_i_60_98 (.ZN(per_dout_mpy[15]), .A(
      multiplier_0_n_60_81), .B1(multiplier_0_n_60_82), .B2(multiplier_0_n_60_7));
  AOI22_X1_LVT multiplier_0_i_60_87 (.ZN(multiplier_0_n_60_73), .A1(
      multiplier_0_n_60_0), .A2(multiplier_0_n_90), .B1(multiplier_0_cycle[1]), 
      .B2(multiplier_0_n_136));
  NOR2_X1_LVT multiplier_0_i_60_88 (.ZN(multiplier_0_n_60_74), .A1(
      multiplier_0_n_60_73), .A2(multiplier_0_n_60_2));
  AND2_X1_LVT multiplier_0_i_60_89 (.ZN(multiplier_0_n_60_75), .A1(
      multiplier_0_n_150), .A2(multiplier_0_op1[14]));
  AND2_X1_LVT multiplier_0_i_19_0 (.ZN(multiplier_0_n_36), .A1(
      multiplier_0_op2_reg[14]), .A2(multiplier_0_n_12));
  NOR4_X1_LVT multiplier_0_i_60_90 (.ZN(multiplier_0_n_60_76), .A1(
      multiplier_0_n_60_74), .A2(multiplier_0_n_60_75), .A3(multiplier_0_n_149), 
      .A4(multiplier_0_n_36));
  AOI22_X1_LVT multiplier_0_i_60_91 (.ZN(multiplier_0_n_60_77), .A1(
      multiplier_0_n_60_0), .A2(multiplier_0_reshi[14]), .B1(
      multiplier_0_cycle[1]), .B2(multiplier_0_reshi_nxt[14]));
  OAI21_X1_LVT multiplier_0_i_60_92 (.ZN(per_dout_mpy[14]), .A(
      multiplier_0_n_60_76), .B1(multiplier_0_n_60_77), .B2(multiplier_0_n_60_7));
  AOI22_X1_LVT multiplier_0_i_60_81 (.ZN(multiplier_0_n_60_68), .A1(
      multiplier_0_n_60_0), .A2(multiplier_0_n_91), .B1(multiplier_0_cycle[1]), 
      .B2(multiplier_0_n_135));
  NOR2_X1_LVT multiplier_0_i_60_82 (.ZN(multiplier_0_n_60_69), .A1(
      multiplier_0_n_60_68), .A2(multiplier_0_n_60_2));
  AND2_X1_LVT multiplier_0_i_60_83 (.ZN(multiplier_0_n_60_70), .A1(
      multiplier_0_n_150), .A2(multiplier_0_op1[13]));
  AND2_X1_LVT multiplier_0_i_18_0 (.ZN(multiplier_0_n_35), .A1(
      multiplier_0_op2_reg[13]), .A2(multiplier_0_n_12));
  NOR4_X1_LVT multiplier_0_i_60_84 (.ZN(multiplier_0_n_60_71), .A1(
      multiplier_0_n_60_69), .A2(multiplier_0_n_60_70), .A3(multiplier_0_n_149), 
      .A4(multiplier_0_n_35));
  AOI22_X1_LVT multiplier_0_i_60_85 (.ZN(multiplier_0_n_60_72), .A1(
      multiplier_0_n_60_0), .A2(multiplier_0_reshi[13]), .B1(
      multiplier_0_cycle[1]), .B2(multiplier_0_reshi_nxt[13]));
  OAI21_X1_LVT multiplier_0_i_60_86 (.ZN(per_dout_mpy[13]), .A(
      multiplier_0_n_60_71), .B1(multiplier_0_n_60_72), .B2(multiplier_0_n_60_7));
  AOI22_X1_LVT multiplier_0_i_60_75 (.ZN(multiplier_0_n_60_63), .A1(
      multiplier_0_n_60_0), .A2(multiplier_0_n_92), .B1(multiplier_0_cycle[1]), 
      .B2(multiplier_0_n_134));
  NOR2_X1_LVT multiplier_0_i_60_76 (.ZN(multiplier_0_n_60_64), .A1(
      multiplier_0_n_60_63), .A2(multiplier_0_n_60_2));
  AND2_X1_LVT multiplier_0_i_60_77 (.ZN(multiplier_0_n_60_65), .A1(
      multiplier_0_n_150), .A2(multiplier_0_op1[12]));
  AND2_X1_LVT multiplier_0_i_17_0 (.ZN(multiplier_0_n_34), .A1(
      multiplier_0_op2_reg[12]), .A2(multiplier_0_n_12));
  NOR4_X1_LVT multiplier_0_i_60_78 (.ZN(multiplier_0_n_60_66), .A1(
      multiplier_0_n_60_64), .A2(multiplier_0_n_60_65), .A3(multiplier_0_n_149), 
      .A4(multiplier_0_n_34));
  AOI22_X1_LVT multiplier_0_i_60_79 (.ZN(multiplier_0_n_60_67), .A1(
      multiplier_0_n_60_0), .A2(multiplier_0_reshi[12]), .B1(
      multiplier_0_cycle[1]), .B2(multiplier_0_reshi_nxt[12]));
  OAI21_X1_LVT multiplier_0_i_60_80 (.ZN(per_dout_mpy[12]), .A(
      multiplier_0_n_60_66), .B1(multiplier_0_n_60_67), .B2(multiplier_0_n_60_7));
  AOI22_X1_LVT multiplier_0_i_60_69 (.ZN(multiplier_0_n_60_58), .A1(
      multiplier_0_n_60_0), .A2(multiplier_0_n_93), .B1(multiplier_0_cycle[1]), 
      .B2(multiplier_0_n_133));
  NOR2_X1_LVT multiplier_0_i_60_70 (.ZN(multiplier_0_n_60_59), .A1(
      multiplier_0_n_60_58), .A2(multiplier_0_n_60_2));
  AND2_X1_LVT multiplier_0_i_60_71 (.ZN(multiplier_0_n_60_60), .A1(
      multiplier_0_n_150), .A2(multiplier_0_op1[11]));
  AND2_X1_LVT multiplier_0_i_16_0 (.ZN(multiplier_0_n_33), .A1(
      multiplier_0_op2_reg[11]), .A2(multiplier_0_n_12));
  NOR4_X1_LVT multiplier_0_i_60_72 (.ZN(multiplier_0_n_60_61), .A1(
      multiplier_0_n_60_59), .A2(multiplier_0_n_60_60), .A3(multiplier_0_n_149), 
      .A4(multiplier_0_n_33));
  AOI22_X1_LVT multiplier_0_i_60_73 (.ZN(multiplier_0_n_60_62), .A1(
      multiplier_0_n_60_0), .A2(multiplier_0_reshi[11]), .B1(
      multiplier_0_cycle[1]), .B2(multiplier_0_reshi_nxt[11]));
  OAI21_X1_LVT multiplier_0_i_60_74 (.ZN(per_dout_mpy[11]), .A(
      multiplier_0_n_60_61), .B1(multiplier_0_n_60_62), .B2(multiplier_0_n_60_7));
  AOI22_X1_LVT multiplier_0_i_60_63 (.ZN(multiplier_0_n_60_53), .A1(
      multiplier_0_n_60_0), .A2(multiplier_0_n_94), .B1(multiplier_0_cycle[1]), 
      .B2(multiplier_0_n_132));
  NOR2_X1_LVT multiplier_0_i_60_64 (.ZN(multiplier_0_n_60_54), .A1(
      multiplier_0_n_60_53), .A2(multiplier_0_n_60_2));
  AND2_X1_LVT multiplier_0_i_60_65 (.ZN(multiplier_0_n_60_55), .A1(
      multiplier_0_n_150), .A2(multiplier_0_op1[10]));
  AND2_X1_LVT multiplier_0_i_15_0 (.ZN(multiplier_0_n_32), .A1(
      multiplier_0_op2_reg[10]), .A2(multiplier_0_n_12));
  NOR4_X1_LVT multiplier_0_i_60_66 (.ZN(multiplier_0_n_60_56), .A1(
      multiplier_0_n_60_54), .A2(multiplier_0_n_60_55), .A3(multiplier_0_n_149), 
      .A4(multiplier_0_n_32));
  AOI22_X1_LVT multiplier_0_i_60_67 (.ZN(multiplier_0_n_60_57), .A1(
      multiplier_0_n_60_0), .A2(multiplier_0_reshi[10]), .B1(
      multiplier_0_cycle[1]), .B2(multiplier_0_reshi_nxt[10]));
  OAI21_X1_LVT multiplier_0_i_60_68 (.ZN(per_dout_mpy[10]), .A(
      multiplier_0_n_60_56), .B1(multiplier_0_n_60_57), .B2(multiplier_0_n_60_7));
  AOI22_X1_LVT multiplier_0_i_60_57 (.ZN(multiplier_0_n_60_48), .A1(
      multiplier_0_n_60_0), .A2(multiplier_0_n_95), .B1(multiplier_0_cycle[1]), 
      .B2(multiplier_0_n_131));
  NOR2_X1_LVT multiplier_0_i_60_58 (.ZN(multiplier_0_n_60_49), .A1(
      multiplier_0_n_60_48), .A2(multiplier_0_n_60_2));
  AND2_X1_LVT multiplier_0_i_60_59 (.ZN(multiplier_0_n_60_50), .A1(
      multiplier_0_n_150), .A2(multiplier_0_op1[9]));
  AND2_X1_LVT multiplier_0_i_14_0 (.ZN(multiplier_0_n_31), .A1(
      multiplier_0_op2_reg[9]), .A2(multiplier_0_n_12));
  NOR4_X1_LVT multiplier_0_i_60_60 (.ZN(multiplier_0_n_60_51), .A1(
      multiplier_0_n_60_49), .A2(multiplier_0_n_60_50), .A3(multiplier_0_n_149), 
      .A4(multiplier_0_n_31));
  AOI22_X1_LVT multiplier_0_i_60_61 (.ZN(multiplier_0_n_60_52), .A1(
      multiplier_0_n_60_0), .A2(multiplier_0_reshi[9]), .B1(
      multiplier_0_cycle[1]), .B2(multiplier_0_reshi_nxt[9]));
  OAI21_X1_LVT multiplier_0_i_60_62 (.ZN(per_dout_mpy[9]), .A(
      multiplier_0_n_60_51), .B1(multiplier_0_n_60_52), .B2(multiplier_0_n_60_7));
  AOI22_X1_LVT multiplier_0_i_60_51 (.ZN(multiplier_0_n_60_43), .A1(
      multiplier_0_n_60_0), .A2(multiplier_0_n_96), .B1(multiplier_0_cycle[1]), 
      .B2(multiplier_0_n_130));
  NOR2_X1_LVT multiplier_0_i_60_52 (.ZN(multiplier_0_n_60_44), .A1(
      multiplier_0_n_60_43), .A2(multiplier_0_n_60_2));
  AND2_X1_LVT multiplier_0_i_60_53 (.ZN(multiplier_0_n_60_45), .A1(
      multiplier_0_n_150), .A2(multiplier_0_op1[8]));
  AND2_X1_LVT multiplier_0_i_13_0 (.ZN(multiplier_0_n_30), .A1(
      multiplier_0_op2_reg[8]), .A2(multiplier_0_n_12));
  NOR4_X1_LVT multiplier_0_i_60_54 (.ZN(multiplier_0_n_60_46), .A1(
      multiplier_0_n_60_44), .A2(multiplier_0_n_60_45), .A3(multiplier_0_n_149), 
      .A4(multiplier_0_n_30));
  AOI22_X1_LVT multiplier_0_i_60_55 (.ZN(multiplier_0_n_60_47), .A1(
      multiplier_0_n_60_0), .A2(multiplier_0_reshi[8]), .B1(
      multiplier_0_cycle[1]), .B2(multiplier_0_reshi_nxt[8]));
  OAI21_X1_LVT multiplier_0_i_60_56 (.ZN(per_dout_mpy[8]), .A(
      multiplier_0_n_60_46), .B1(multiplier_0_n_60_47), .B2(multiplier_0_n_60_7));
  AOI22_X1_LVT multiplier_0_i_60_45 (.ZN(multiplier_0_n_60_38), .A1(
      multiplier_0_n_60_0), .A2(multiplier_0_n_97), .B1(multiplier_0_cycle[1]), 
      .B2(multiplier_0_n_129));
  NOR2_X1_LVT multiplier_0_i_60_46 (.ZN(multiplier_0_n_60_39), .A1(
      multiplier_0_n_60_38), .A2(multiplier_0_n_60_2));
  AND2_X1_LVT multiplier_0_i_60_47 (.ZN(multiplier_0_n_60_40), .A1(
      multiplier_0_n_150), .A2(multiplier_0_op1[7]));
  AND2_X1_LVT multiplier_0_i_12_7 (.ZN(multiplier_0_n_29), .A1(multiplier_0_n_12), 
      .A2(multiplier_0_op2_reg[7]));
  NOR4_X1_LVT multiplier_0_i_60_48 (.ZN(multiplier_0_n_60_41), .A1(
      multiplier_0_n_60_39), .A2(multiplier_0_n_60_40), .A3(multiplier_0_n_149), 
      .A4(multiplier_0_n_29));
  AOI22_X1_LVT multiplier_0_i_60_49 (.ZN(multiplier_0_n_60_42), .A1(
      multiplier_0_n_60_0), .A2(multiplier_0_reshi[7]), .B1(
      multiplier_0_cycle[1]), .B2(multiplier_0_reshi_nxt[7]));
  OAI21_X1_LVT multiplier_0_i_60_50 (.ZN(per_dout_mpy[7]), .A(
      multiplier_0_n_60_41), .B1(multiplier_0_n_60_42), .B2(multiplier_0_n_60_7));
  AOI22_X1_LVT multiplier_0_i_60_39 (.ZN(multiplier_0_n_60_33), .A1(
      multiplier_0_n_60_0), .A2(multiplier_0_n_98), .B1(multiplier_0_cycle[1]), 
      .B2(multiplier_0_n_128));
  NOR2_X1_LVT multiplier_0_i_60_40 (.ZN(multiplier_0_n_60_34), .A1(
      multiplier_0_n_60_33), .A2(multiplier_0_n_60_2));
  AND2_X1_LVT multiplier_0_i_60_41 (.ZN(multiplier_0_n_60_35), .A1(
      multiplier_0_n_150), .A2(multiplier_0_op1[6]));
  AND2_X1_LVT multiplier_0_i_12_6 (.ZN(multiplier_0_n_28), .A1(multiplier_0_n_12), 
      .A2(multiplier_0_op2_reg[6]));
  NOR4_X1_LVT multiplier_0_i_60_42 (.ZN(multiplier_0_n_60_36), .A1(
      multiplier_0_n_60_34), .A2(multiplier_0_n_60_35), .A3(multiplier_0_n_149), 
      .A4(multiplier_0_n_28));
  AOI22_X1_LVT multiplier_0_i_60_43 (.ZN(multiplier_0_n_60_37), .A1(
      multiplier_0_n_60_0), .A2(multiplier_0_reshi[6]), .B1(
      multiplier_0_cycle[1]), .B2(multiplier_0_reshi_nxt[6]));
  OAI21_X1_LVT multiplier_0_i_60_44 (.ZN(per_dout_mpy[6]), .A(
      multiplier_0_n_60_36), .B1(multiplier_0_n_60_37), .B2(multiplier_0_n_60_7));
  AOI22_X1_LVT multiplier_0_i_60_33 (.ZN(multiplier_0_n_60_28), .A1(
      multiplier_0_n_60_0), .A2(multiplier_0_n_99), .B1(multiplier_0_cycle[1]), 
      .B2(multiplier_0_n_127));
  NOR2_X1_LVT multiplier_0_i_60_34 (.ZN(multiplier_0_n_60_29), .A1(
      multiplier_0_n_60_28), .A2(multiplier_0_n_60_2));
  AND2_X1_LVT multiplier_0_i_60_35 (.ZN(multiplier_0_n_60_30), .A1(
      multiplier_0_n_150), .A2(multiplier_0_op1[5]));
  AND2_X1_LVT multiplier_0_i_12_5 (.ZN(multiplier_0_n_27), .A1(multiplier_0_n_12), 
      .A2(multiplier_0_op2_reg[5]));
  NOR4_X1_LVT multiplier_0_i_60_36 (.ZN(multiplier_0_n_60_31), .A1(
      multiplier_0_n_60_29), .A2(multiplier_0_n_60_30), .A3(multiplier_0_n_149), 
      .A4(multiplier_0_n_27));
  AOI22_X1_LVT multiplier_0_i_60_37 (.ZN(multiplier_0_n_60_32), .A1(
      multiplier_0_n_60_0), .A2(multiplier_0_reshi[5]), .B1(
      multiplier_0_cycle[1]), .B2(multiplier_0_reshi_nxt[5]));
  OAI21_X1_LVT multiplier_0_i_60_38 (.ZN(per_dout_mpy[5]), .A(
      multiplier_0_n_60_31), .B1(multiplier_0_n_60_32), .B2(multiplier_0_n_60_7));
  AOI22_X1_LVT multiplier_0_i_60_27 (.ZN(multiplier_0_n_60_23), .A1(
      multiplier_0_n_60_0), .A2(multiplier_0_n_100), .B1(multiplier_0_cycle[1]), 
      .B2(multiplier_0_n_126));
  NOR2_X1_LVT multiplier_0_i_60_28 (.ZN(multiplier_0_n_60_24), .A1(
      multiplier_0_n_60_23), .A2(multiplier_0_n_60_2));
  AND2_X1_LVT multiplier_0_i_60_29 (.ZN(multiplier_0_n_60_25), .A1(
      multiplier_0_n_150), .A2(multiplier_0_op1[4]));
  AND2_X1_LVT multiplier_0_i_12_4 (.ZN(multiplier_0_n_26), .A1(multiplier_0_n_12), 
      .A2(multiplier_0_op2_reg[4]));
  NOR4_X1_LVT multiplier_0_i_60_30 (.ZN(multiplier_0_n_60_26), .A1(
      multiplier_0_n_60_24), .A2(multiplier_0_n_60_25), .A3(multiplier_0_n_149), 
      .A4(multiplier_0_n_26));
  AOI22_X1_LVT multiplier_0_i_60_31 (.ZN(multiplier_0_n_60_27), .A1(
      multiplier_0_n_60_0), .A2(multiplier_0_reshi[4]), .B1(
      multiplier_0_cycle[1]), .B2(multiplier_0_reshi_nxt[4]));
  OAI21_X1_LVT multiplier_0_i_60_32 (.ZN(per_dout_mpy[4]), .A(
      multiplier_0_n_60_26), .B1(multiplier_0_n_60_27), .B2(multiplier_0_n_60_7));
  AOI22_X1_LVT multiplier_0_i_60_21 (.ZN(multiplier_0_n_60_18), .A1(
      multiplier_0_n_60_0), .A2(multiplier_0_n_101), .B1(multiplier_0_cycle[1]), 
      .B2(multiplier_0_n_125));
  NOR2_X1_LVT multiplier_0_i_60_22 (.ZN(multiplier_0_n_60_19), .A1(
      multiplier_0_n_60_18), .A2(multiplier_0_n_60_2));
  AND2_X1_LVT multiplier_0_i_60_23 (.ZN(multiplier_0_n_60_20), .A1(
      multiplier_0_n_150), .A2(multiplier_0_op1[3]));
  AND2_X1_LVT multiplier_0_i_12_3 (.ZN(multiplier_0_n_25), .A1(multiplier_0_n_12), 
      .A2(multiplier_0_op2_reg[3]));
  NOR4_X1_LVT multiplier_0_i_60_24 (.ZN(multiplier_0_n_60_21), .A1(
      multiplier_0_n_60_19), .A2(multiplier_0_n_60_20), .A3(multiplier_0_n_149), 
      .A4(multiplier_0_n_25));
  AOI22_X1_LVT multiplier_0_i_60_25 (.ZN(multiplier_0_n_60_22), .A1(
      multiplier_0_n_60_0), .A2(multiplier_0_reshi[3]), .B1(
      multiplier_0_cycle[1]), .B2(multiplier_0_reshi_nxt[3]));
  OAI21_X1_LVT multiplier_0_i_60_26 (.ZN(per_dout_mpy[3]), .A(
      multiplier_0_n_60_21), .B1(multiplier_0_n_60_22), .B2(multiplier_0_n_60_7));
  AOI22_X1_LVT multiplier_0_i_60_15 (.ZN(multiplier_0_n_60_13), .A1(
      multiplier_0_n_60_0), .A2(multiplier_0_n_102), .B1(multiplier_0_cycle[1]), 
      .B2(multiplier_0_n_124));
  NOR2_X1_LVT multiplier_0_i_60_16 (.ZN(multiplier_0_n_60_14), .A1(
      multiplier_0_n_60_13), .A2(multiplier_0_n_60_2));
  AND2_X1_LVT multiplier_0_i_60_17 (.ZN(multiplier_0_n_60_15), .A1(
      multiplier_0_n_150), .A2(multiplier_0_op1[2]));
  AND2_X1_LVT multiplier_0_i_12_2 (.ZN(multiplier_0_n_24), .A1(multiplier_0_n_12), 
      .A2(multiplier_0_op2_reg[2]));
  NOR4_X1_LVT multiplier_0_i_60_18 (.ZN(multiplier_0_n_60_16), .A1(
      multiplier_0_n_60_14), .A2(multiplier_0_n_60_15), .A3(multiplier_0_n_149), 
      .A4(multiplier_0_n_24));
  AOI22_X1_LVT multiplier_0_i_60_19 (.ZN(multiplier_0_n_60_17), .A1(
      multiplier_0_n_60_0), .A2(multiplier_0_reshi[2]), .B1(
      multiplier_0_cycle[1]), .B2(multiplier_0_reshi_nxt[2]));
  OAI21_X1_LVT multiplier_0_i_60_20 (.ZN(per_dout_mpy[2]), .A(
      multiplier_0_n_60_16), .B1(multiplier_0_n_60_17), .B2(multiplier_0_n_60_7));
  AOI22_X1_LVT multiplier_0_i_60_9 (.ZN(multiplier_0_n_60_8), .A1(
      multiplier_0_n_60_0), .A2(multiplier_0_n_103), .B1(multiplier_0_cycle[1]), 
      .B2(multiplier_0_n_123));
  NOR2_X1_LVT multiplier_0_i_60_10 (.ZN(multiplier_0_n_60_9), .A1(
      multiplier_0_n_60_8), .A2(multiplier_0_n_60_2));
  AND2_X1_LVT multiplier_0_i_60_11 (.ZN(multiplier_0_n_60_10), .A1(
      multiplier_0_n_150), .A2(multiplier_0_op1[1]));
  INV_X1_LVT multiplier_0_i_55_0 (.ZN(multiplier_0_n_55_0), .A(
      multiplier_0_cycle[1]));
  AOI22_X1_LVT multiplier_0_i_55_3 (.ZN(multiplier_0_n_55_2), .A1(
      multiplier_0_n_55_0), .A2(multiplier_0_sumext_s[1]), .B1(
      multiplier_0_cycle[1]), .B2(multiplier_0_sumext_s_nxt[1]));
  INV_X1_LVT multiplier_0_i_55_4 (.ZN(multiplier_0_n_145), .A(
      multiplier_0_n_55_2));
  AND2_X1_LVT multiplier_0_i_56_1 (.ZN(multiplier_0_n_147), .A1(
      multiplier_0_reg_rd15), .A2(multiplier_0_n_145));
  AND2_X1_LVT multiplier_0_i_12_1 (.ZN(multiplier_0_n_23), .A1(multiplier_0_n_12), 
      .A2(multiplier_0_op2_reg[1]));
  NOR4_X1_LVT multiplier_0_i_60_12 (.ZN(multiplier_0_n_60_11), .A1(
      multiplier_0_n_60_9), .A2(multiplier_0_n_60_10), .A3(multiplier_0_n_147), 
      .A4(multiplier_0_n_23));
  AOI22_X1_LVT multiplier_0_i_60_13 (.ZN(multiplier_0_n_60_12), .A1(
      multiplier_0_n_60_0), .A2(multiplier_0_reshi[1]), .B1(
      multiplier_0_cycle[1]), .B2(multiplier_0_reshi_nxt[1]));
  OAI21_X1_LVT multiplier_0_i_60_14 (.ZN(per_dout_mpy[1]), .A(
      multiplier_0_n_60_11), .B1(multiplier_0_n_60_12), .B2(multiplier_0_n_60_7));
  AOI22_X1_LVT multiplier_0_i_60_1 (.ZN(multiplier_0_n_60_1), .A1(
      multiplier_0_n_60_0), .A2(multiplier_0_n_104), .B1(multiplier_0_cycle[1]), 
      .B2(multiplier_0_n_122));
  NOR2_X1_LVT multiplier_0_i_60_3 (.ZN(multiplier_0_n_60_3), .A1(
      multiplier_0_n_60_1), .A2(multiplier_0_n_60_2));
  AND2_X1_LVT multiplier_0_i_60_4 (.ZN(multiplier_0_n_60_4), .A1(
      multiplier_0_op1[0]), .A2(multiplier_0_n_150));
  OR2_X1_LVT multiplier_0_i_49_0 (.ZN(multiplier_0_n_139), .A1(
      multiplier_0_n_138), .A2(multiplier_0_sumext_s[0]));
  INV_X1_LVT multiplier_0_i_50_1 (.ZN(multiplier_0_n_50_1), .A(
      multiplier_0_n_139));
  OAI21_X1_LVT multiplier_0_i_50_2 (.ZN(multiplier_0_sumext_s_nxt[0]), .A(
      multiplier_0_n_50_0), .B1(multiplier_0_n_50_1), .B2(multiplier_0_sign_sel));
  AND2_X1_LVT multiplier_0_i_52_1 (.ZN(multiplier_0_n_141), .A1(
      multiplier_0_n_52_0), .A2(multiplier_0_sumext_s_nxt[0]));
  DFFR_X1_LVT \multiplier_0_sumext_s_reg[0] (.Q(multiplier_0_sumext_s[0]), .QN(), 
      .CK(multiplier_0_n_140), .D(multiplier_0_n_141), .RN(multiplier_0_n_38));
  AOI22_X1_LVT multiplier_0_i_55_1 (.ZN(multiplier_0_n_55_1), .A1(
      multiplier_0_n_55_0), .A2(multiplier_0_sumext_s[0]), .B1(
      multiplier_0_sumext_s_nxt[0]), .B2(multiplier_0_cycle[1]));
  INV_X1_LVT multiplier_0_i_55_2 (.ZN(multiplier_0_n_144), .A(
      multiplier_0_n_55_1));
  AND2_X1_LVT multiplier_0_i_56_0 (.ZN(multiplier_0_n_146), .A1(
      multiplier_0_n_144), .A2(multiplier_0_reg_rd15));
  AND2_X1_LVT multiplier_0_i_12_0 (.ZN(multiplier_0_n_22), .A1(
      multiplier_0_op2_reg[0]), .A2(multiplier_0_n_12));
  NOR4_X1_LVT multiplier_0_i_60_5 (.ZN(multiplier_0_n_60_5), .A1(
      multiplier_0_n_60_3), .A2(multiplier_0_n_60_4), .A3(multiplier_0_n_146), 
      .A4(multiplier_0_n_22));
  AOI22_X1_LVT multiplier_0_i_60_6 (.ZN(multiplier_0_n_60_6), .A1(
      multiplier_0_n_60_0), .A2(multiplier_0_reshi[0]), .B1(
      multiplier_0_reshi_nxt[0]), .B2(multiplier_0_cycle[1]));
  OAI21_X1_LVT multiplier_0_i_60_8 (.ZN(per_dout_mpy[0]), .A(multiplier_0_n_60_5), 
      .B1(multiplier_0_n_60_6), .B2(multiplier_0_n_60_7));
  OR4_X1_LVT i_0_0_30 (.ZN(n_0_0_15), .A1(per_dout_mpy[15]), .A2(
      per_dout_wdog[15]), .A3(per_dout_sfr[15]), .A4(per_dout_clk[15]));
  OR2_X1_LVT i_0_0_31 (.ZN(per_dout_or[15]), .A1(n_0_0_15), .A2(per_dout[15]));
  OR4_X1_LVT i_0_0_28 (.ZN(n_0_0_14), .A1(per_dout_mpy[14]), .A2(
      per_dout_wdog[14]), .A3(per_dout_sfr[14]), .A4(per_dout_clk[14]));
  OR2_X1_LVT i_0_0_29 (.ZN(per_dout_or[14]), .A1(n_0_0_14), .A2(per_dout[14]));
  OR4_X1_LVT i_0_0_26 (.ZN(n_0_0_13), .A1(per_dout_mpy[13]), .A2(
      per_dout_wdog[13]), .A3(per_dout_sfr[13]), .A4(per_dout_clk[13]));
  OR2_X1_LVT i_0_0_27 (.ZN(per_dout_or[13]), .A1(n_0_0_13), .A2(per_dout[13]));
  OR4_X1_LVT i_0_0_24 (.ZN(n_0_0_12), .A1(per_dout_mpy[12]), .A2(
      per_dout_wdog[12]), .A3(per_dout_sfr[12]), .A4(per_dout_clk[12]));
  OR2_X1_LVT i_0_0_25 (.ZN(per_dout_or[12]), .A1(n_0_0_12), .A2(per_dout[12]));
  OR4_X1_LVT i_0_0_22 (.ZN(n_0_0_11), .A1(per_dout_mpy[11]), .A2(
      per_dout_wdog[11]), .A3(per_dout_sfr[11]), .A4(per_dout_clk[11]));
  OR2_X1_LVT i_0_0_23 (.ZN(per_dout_or[11]), .A1(n_0_0_11), .A2(per_dout[11]));
  OR4_X1_LVT i_0_0_20 (.ZN(n_0_0_10), .A1(per_dout_mpy[10]), .A2(
      per_dout_wdog[10]), .A3(per_dout_sfr[10]), .A4(per_dout_clk[10]));
  OR2_X1_LVT i_0_0_21 (.ZN(per_dout_or[10]), .A1(n_0_0_10), .A2(per_dout[10]));
  OR4_X1_LVT i_0_0_18 (.ZN(n_0_0_9), .A1(per_dout_mpy[9]), .A2(per_dout_wdog[9]), 
      .A3(per_dout_sfr[9]), .A4(per_dout_clk[9]));
  OR2_X1_LVT i_0_0_19 (.ZN(per_dout_or[9]), .A1(n_0_0_9), .A2(per_dout[9]));
  OR4_X1_LVT i_0_0_16 (.ZN(n_0_0_8), .A1(per_dout_mpy[8]), .A2(per_dout_wdog[8]), 
      .A3(per_dout_sfr[8]), .A4(per_dout_clk[8]));
  OR2_X1_LVT i_0_0_17 (.ZN(per_dout_or[8]), .A1(n_0_0_8), .A2(per_dout[8]));
  OR4_X1_LVT i_0_0_14 (.ZN(n_0_0_7), .A1(per_dout_mpy[7]), .A2(per_dout_wdog[7]), 
      .A3(per_dout_sfr[7]), .A4(per_dout_clk[7]));
  OR2_X1_LVT i_0_0_15 (.ZN(per_dout_or[7]), .A1(n_0_0_7), .A2(per_dout[7]));
  OR4_X1_LVT i_0_0_12 (.ZN(n_0_0_6), .A1(per_dout_mpy[6]), .A2(per_dout_wdog[6]), 
      .A3(per_dout_sfr[6]), .A4(per_dout_clk[6]));
  OR2_X1_LVT i_0_0_13 (.ZN(per_dout_or[6]), .A1(n_0_0_6), .A2(per_dout[6]));
  OR4_X1_LVT i_0_0_10 (.ZN(n_0_0_5), .A1(per_dout_mpy[5]), .A2(per_dout_wdog[5]), 
      .A3(per_dout_sfr[5]), .A4(per_dout_clk[5]));
  OR2_X1_LVT i_0_0_11 (.ZN(per_dout_or[5]), .A1(n_0_0_5), .A2(per_dout[5]));
  OR4_X1_LVT i_0_0_8 (.ZN(n_0_0_4), .A1(per_dout_mpy[4]), .A2(per_dout_wdog[4]), 
      .A3(per_dout_sfr[4]), .A4(per_dout_clk[4]));
  OR2_X1_LVT i_0_0_9 (.ZN(per_dout_or[4]), .A1(n_0_0_4), .A2(per_dout[4]));
  OR4_X1_LVT i_0_0_6 (.ZN(n_0_0_3), .A1(per_dout_mpy[3]), .A2(per_dout_wdog[3]), 
      .A3(per_dout_sfr[3]), .A4(per_dout_clk[3]));
  OR2_X1_LVT i_0_0_7 (.ZN(per_dout_or[3]), .A1(n_0_0_3), .A2(per_dout[3]));
  OR4_X1_LVT i_0_0_4 (.ZN(n_0_0_2), .A1(per_dout_mpy[2]), .A2(per_dout_wdog[2]), 
      .A3(per_dout_sfr[2]), .A4(per_dout_clk[2]));
  OR2_X1_LVT i_0_0_5 (.ZN(per_dout_or[2]), .A1(n_0_0_2), .A2(per_dout[2]));
  OR4_X1_LVT i_0_0_2 (.ZN(n_0_0_1), .A1(per_dout_mpy[1]), .A2(per_dout_wdog[1]), 
      .A3(per_dout_sfr[1]), .A4(per_dout_clk[1]));
  OR2_X1_LVT i_0_0_3 (.ZN(per_dout_or[1]), .A1(n_0_0_1), .A2(per_dout[1]));
  OR4_X1_LVT i_0_0_0 (.ZN(n_0_0_0), .A1(per_dout_mpy[0]), .A2(per_dout_wdog[0]), 
      .A3(per_dout_sfr[0]), .A4(per_dout_clk[0]));
  OR2_X1_LVT i_0_0_1 (.ZN(per_dout_or[0]), .A1(n_0_0_0), .A2(per_dout[0]));
  AOI21_X1_LVT mem_backbone_0_i_0_0 (.ZN(mem_backbone_0_n_0_0), .A(dbg_halt_cmd), 
      .B1(dma_en), .B2(dma_priority));
  INV_X1_LVT mem_backbone_0_i_0_1 (.ZN(cpu_halt_cmd), .A(mem_backbone_0_n_0_0));
  OR2_X1_LVT mem_backbone_0_i_4_0 (.ZN(mem_backbone_0_ext_mem_en), .A1(
      dbg_mem_en), .A2(dma_en));
  AND4_X1_LVT mem_backbone_0_i_8_0 (.ZN(mem_backbone_0_n_8_0), .A1(n_12), .A2(
      n_13), .A3(n_14), .A4(fe_mb_en));
  AND2_X1_LVT mem_backbone_0_i_8_1 (.ZN(mem_backbone_0_fe_pmem_en), .A1(
      mem_backbone_0_n_8_0), .A2(n_11));
  INV_X1_LVT mem_backbone_0_i_9_0 (.ZN(mem_backbone_0_n_0), .A(
      mem_backbone_0_fe_pmem_en));
  INV_X1_LVT mem_backbone_0_i_2_0 (.ZN(mem_backbone_0_n_2_0), .A(dbg_mem_en));
  AOI22_X1_LVT mem_backbone_0_i_2_23 (.ZN(mem_backbone_0_n_2_12), .A1(
      mem_backbone_0_n_2_0), .A2(dma_addr[11]), .B1(dbg_mem_en), .B2(
      dbg_mem_addr[12]));
  INV_X1_LVT mem_backbone_0_i_2_24 (.ZN(mem_backbone_0_ext_mem_addr[11]), .A(
      mem_backbone_0_n_2_12));
  AOI22_X1_LVT mem_backbone_0_i_2_25 (.ZN(mem_backbone_0_n_2_13), .A1(
      mem_backbone_0_n_2_0), .A2(dma_addr[12]), .B1(dbg_mem_en), .B2(
      dbg_mem_addr[13]));
  INV_X1_LVT mem_backbone_0_i_2_26 (.ZN(mem_backbone_0_ext_mem_addr[12]), .A(
      mem_backbone_0_n_2_13));
  AOI22_X1_LVT mem_backbone_0_i_2_27 (.ZN(mem_backbone_0_n_2_14), .A1(
      mem_backbone_0_n_2_0), .A2(dma_addr[13]), .B1(dbg_mem_en), .B2(
      dbg_mem_addr[14]));
  INV_X1_LVT mem_backbone_0_i_2_28 (.ZN(mem_backbone_0_ext_mem_addr[13]), .A(
      mem_backbone_0_n_2_14));
  AOI22_X1_LVT mem_backbone_0_i_2_29 (.ZN(mem_backbone_0_n_2_15), .A1(
      mem_backbone_0_n_2_0), .A2(dma_addr[14]), .B1(dbg_mem_en), .B2(
      dbg_mem_addr[15]));
  INV_X1_LVT mem_backbone_0_i_2_30 (.ZN(mem_backbone_0_ext_mem_addr[14]), .A(
      mem_backbone_0_n_2_15));
  AND4_X1_LVT mem_backbone_0_i_7_0 (.ZN(mem_backbone_0_ext_pmem_sel), .A1(
      mem_backbone_0_ext_mem_addr[11]), .A2(mem_backbone_0_ext_mem_addr[12]), 
      .A3(mem_backbone_0_ext_mem_addr[13]), .A4(mem_backbone_0_ext_mem_addr[14]));
  NAND3_X1_LVT mem_backbone_0_i_12_0 (.ZN(mem_backbone_0_n_12_0), .A1(
      mem_backbone_0_ext_mem_en), .A2(mem_backbone_0_n_0), .A3(
      mem_backbone_0_ext_pmem_sel));
  NOR2_X1_LVT mem_backbone_0_i_10_0 (.ZN(mem_backbone_0_n_1), .A1(eu_mb_wr[0]), 
      .A2(eu_mb_wr[1]));
  NAND4_X1_LVT mem_backbone_0_i_11_0 (.ZN(mem_backbone_0_n_11_0), .A1(eu_mab[14]), 
      .A2(eu_mab[15]), .A3(eu_mb_en), .A4(mem_backbone_0_n_1));
  NAND2_X1_LVT mem_backbone_0_i_11_1 (.ZN(mem_backbone_0_n_11_1), .A1(eu_mab[12]), 
      .A2(eu_mab[13]));
  NOR2_X1_LVT mem_backbone_0_i_11_2 (.ZN(mem_backbone_0_eu_pmem_en), .A1(
      mem_backbone_0_n_11_0), .A2(mem_backbone_0_n_11_1));
  NOR2_X1_LVT mem_backbone_0_i_12_1 (.ZN(mem_backbone_0_ext_pmem_en), .A1(
      mem_backbone_0_n_12_0), .A2(mem_backbone_0_eu_pmem_en));
  INV_X1_LVT mem_backbone_0_i_13_0 (.ZN(mem_backbone_0_n_2), .A(puc_rst));
  DFFR_X1_LVT \mem_backbone_0_ext_mem_din_sel_reg[1] (.Q(
      mem_backbone_0_ext_mem_din_sel[1]), .QN(), .CK(mclk), .D(
      mem_backbone_0_ext_pmem_en), .RN(mem_backbone_0_n_2));
  OR4_X1_LVT mem_backbone_0_i_3_0 (.ZN(mem_backbone_0_n_3_0), .A1(
      mem_backbone_0_ext_mem_addr[11]), .A2(mem_backbone_0_ext_mem_addr[12]), 
      .A3(mem_backbone_0_ext_mem_addr[13]), .A4(mem_backbone_0_ext_mem_addr[14]));
  AOI22_X1_LVT mem_backbone_0_i_2_17 (.ZN(mem_backbone_0_n_2_9), .A1(
      mem_backbone_0_n_2_0), .A2(dma_addr[8]), .B1(dbg_mem_en), .B2(
      dbg_mem_addr[9]));
  INV_X1_LVT mem_backbone_0_i_2_18 (.ZN(mem_backbone_0_ext_mem_addr[8]), .A(
      mem_backbone_0_n_2_9));
  AOI22_X1_LVT mem_backbone_0_i_2_19 (.ZN(mem_backbone_0_n_2_10), .A1(
      mem_backbone_0_n_2_0), .A2(dma_addr[9]), .B1(dbg_mem_en), .B2(
      dbg_mem_addr[10]));
  INV_X1_LVT mem_backbone_0_i_2_20 (.ZN(mem_backbone_0_ext_mem_addr[9]), .A(
      mem_backbone_0_n_2_10));
  AOI22_X1_LVT mem_backbone_0_i_2_21 (.ZN(mem_backbone_0_n_2_11), .A1(
      mem_backbone_0_n_2_0), .A2(dma_addr[10]), .B1(dbg_mem_en), .B2(
      dbg_mem_addr[11]));
  INV_X1_LVT mem_backbone_0_i_2_22 (.ZN(mem_backbone_0_ext_mem_addr[10]), .A(
      mem_backbone_0_n_2_11));
  NOR4_X1_LVT mem_backbone_0_i_3_1 (.ZN(mem_backbone_0_ext_per_sel), .A1(
      mem_backbone_0_n_3_0), .A2(mem_backbone_0_ext_mem_addr[8]), .A3(
      mem_backbone_0_ext_mem_addr[9]), .A4(mem_backbone_0_ext_mem_addr[10]));
  NAND2_X1_LVT mem_backbone_0_i_6_0 (.ZN(mem_backbone_0_n_6_0), .A1(
      mem_backbone_0_ext_mem_en), .A2(mem_backbone_0_ext_per_sel));
  INV_X1_LVT mem_backbone_0_i_5_0 (.ZN(mem_backbone_0_n_5_0), .A(eu_mb_en));
  NOR4_X1_LVT mem_backbone_0_i_5_1 (.ZN(mem_backbone_0_n_5_1), .A1(
      mem_backbone_0_n_5_0), .A2(eu_mab[13]), .A3(eu_mab[14]), .A4(eu_mab[15]));
  NOR4_X1_LVT mem_backbone_0_i_5_2 (.ZN(mem_backbone_0_n_5_2), .A1(eu_mab[9]), 
      .A2(eu_mab[10]), .A3(eu_mab[11]), .A4(eu_mab[12]));
  AND2_X1_LVT mem_backbone_0_i_5_3 (.ZN(mem_backbone_0_eu_per_en), .A1(
      mem_backbone_0_n_5_1), .A2(mem_backbone_0_n_5_2));
  NOR2_X1_LVT mem_backbone_0_i_6_1 (.ZN(mem_backbone_0_ext_per_en), .A1(
      mem_backbone_0_n_6_0), .A2(mem_backbone_0_eu_per_en));
  DFFR_X1_LVT \mem_backbone_0_ext_mem_din_sel_reg[0] (.Q(
      mem_backbone_0_ext_mem_din_sel[0]), .QN(), .CK(mclk), .D(
      mem_backbone_0_ext_per_en), .RN(mem_backbone_0_n_2));
  INV_X1_LVT mem_backbone_0_i_15_1 (.ZN(mem_backbone_0_n_15_0), .A(
      mem_backbone_0_ext_mem_din_sel[0]));
  NOR2_X1_LVT mem_backbone_0_i_15_2 (.ZN(mem_backbone_0_n_4), .A1(
      mem_backbone_0_n_15_0), .A2(mem_backbone_0_ext_mem_din_sel[1]));
  DFFR_X1_LVT \mem_backbone_0_per_dout_val_reg[15] (.Q(
      mem_backbone_0_per_dout_val[15]), .QN(), .CK(mclk), .D(per_dout_or[15]), 
      .RN(mem_backbone_0_n_2));
  NOR2_X1_LVT mem_backbone_0_i_15_0 (.ZN(mem_backbone_0_n_3), .A1(
      mem_backbone_0_ext_mem_din_sel[0]), .A2(mem_backbone_0_ext_mem_din_sel[1]));
  AOI222_X1_LVT mem_backbone_0_i_16_30 (.ZN(mem_backbone_0_n_16_15), .A1(
      mem_backbone_0_ext_mem_din_sel[1]), .A2(pmem_dout[15]), .B1(
      mem_backbone_0_n_4), .B2(mem_backbone_0_per_dout_val[15]), .C1(
      mem_backbone_0_n_3), .C2(dmem_dout[15]));
  INV_X1_LVT mem_backbone_0_i_16_31 (.ZN(dbg_mem_din[15]), .A(
      mem_backbone_0_n_16_15));
  DFFR_X1_LVT \mem_backbone_0_per_dout_val_reg[14] (.Q(
      mem_backbone_0_per_dout_val[14]), .QN(), .CK(mclk), .D(per_dout_or[14]), 
      .RN(mem_backbone_0_n_2));
  AOI222_X1_LVT mem_backbone_0_i_16_28 (.ZN(mem_backbone_0_n_16_14), .A1(
      mem_backbone_0_ext_mem_din_sel[1]), .A2(pmem_dout[14]), .B1(
      mem_backbone_0_n_4), .B2(mem_backbone_0_per_dout_val[14]), .C1(
      mem_backbone_0_n_3), .C2(dmem_dout[14]));
  INV_X1_LVT mem_backbone_0_i_16_29 (.ZN(dbg_mem_din[14]), .A(
      mem_backbone_0_n_16_14));
  DFFR_X1_LVT \mem_backbone_0_per_dout_val_reg[13] (.Q(
      mem_backbone_0_per_dout_val[13]), .QN(), .CK(mclk), .D(per_dout_or[13]), 
      .RN(mem_backbone_0_n_2));
  AOI222_X1_LVT mem_backbone_0_i_16_26 (.ZN(mem_backbone_0_n_16_13), .A1(
      mem_backbone_0_ext_mem_din_sel[1]), .A2(pmem_dout[13]), .B1(
      mem_backbone_0_n_4), .B2(mem_backbone_0_per_dout_val[13]), .C1(
      mem_backbone_0_n_3), .C2(dmem_dout[13]));
  INV_X1_LVT mem_backbone_0_i_16_27 (.ZN(dbg_mem_din[13]), .A(
      mem_backbone_0_n_16_13));
  DFFR_X1_LVT \mem_backbone_0_per_dout_val_reg[12] (.Q(
      mem_backbone_0_per_dout_val[12]), .QN(), .CK(mclk), .D(per_dout_or[12]), 
      .RN(mem_backbone_0_n_2));
  AOI222_X1_LVT mem_backbone_0_i_16_24 (.ZN(mem_backbone_0_n_16_12), .A1(
      mem_backbone_0_ext_mem_din_sel[1]), .A2(pmem_dout[12]), .B1(
      mem_backbone_0_n_4), .B2(mem_backbone_0_per_dout_val[12]), .C1(
      mem_backbone_0_n_3), .C2(dmem_dout[12]));
  INV_X1_LVT mem_backbone_0_i_16_25 (.ZN(dbg_mem_din[12]), .A(
      mem_backbone_0_n_16_12));
  DFFR_X1_LVT \mem_backbone_0_per_dout_val_reg[11] (.Q(
      mem_backbone_0_per_dout_val[11]), .QN(), .CK(mclk), .D(per_dout_or[11]), 
      .RN(mem_backbone_0_n_2));
  AOI222_X1_LVT mem_backbone_0_i_16_22 (.ZN(mem_backbone_0_n_16_11), .A1(
      mem_backbone_0_ext_mem_din_sel[1]), .A2(pmem_dout[11]), .B1(
      mem_backbone_0_n_4), .B2(mem_backbone_0_per_dout_val[11]), .C1(
      mem_backbone_0_n_3), .C2(dmem_dout[11]));
  INV_X1_LVT mem_backbone_0_i_16_23 (.ZN(dbg_mem_din[11]), .A(
      mem_backbone_0_n_16_11));
  DFFR_X1_LVT \mem_backbone_0_per_dout_val_reg[10] (.Q(
      mem_backbone_0_per_dout_val[10]), .QN(), .CK(mclk), .D(per_dout_or[10]), 
      .RN(mem_backbone_0_n_2));
  AOI222_X1_LVT mem_backbone_0_i_16_20 (.ZN(mem_backbone_0_n_16_10), .A1(
      mem_backbone_0_ext_mem_din_sel[1]), .A2(pmem_dout[10]), .B1(
      mem_backbone_0_n_4), .B2(mem_backbone_0_per_dout_val[10]), .C1(
      mem_backbone_0_n_3), .C2(dmem_dout[10]));
  INV_X1_LVT mem_backbone_0_i_16_21 (.ZN(dbg_mem_din[10]), .A(
      mem_backbone_0_n_16_10));
  DFFR_X1_LVT \mem_backbone_0_per_dout_val_reg[9] (.Q(
      mem_backbone_0_per_dout_val[9]), .QN(), .CK(mclk), .D(per_dout_or[9]), .RN(
      mem_backbone_0_n_2));
  AOI222_X1_LVT mem_backbone_0_i_16_18 (.ZN(mem_backbone_0_n_16_9), .A1(
      mem_backbone_0_ext_mem_din_sel[1]), .A2(pmem_dout[9]), .B1(
      mem_backbone_0_n_4), .B2(mem_backbone_0_per_dout_val[9]), .C1(
      mem_backbone_0_n_3), .C2(dmem_dout[9]));
  INV_X1_LVT mem_backbone_0_i_16_19 (.ZN(dbg_mem_din[9]), .A(
      mem_backbone_0_n_16_9));
  DFFR_X1_LVT \mem_backbone_0_per_dout_val_reg[8] (.Q(
      mem_backbone_0_per_dout_val[8]), .QN(), .CK(mclk), .D(per_dout_or[8]), .RN(
      mem_backbone_0_n_2));
  AOI222_X1_LVT mem_backbone_0_i_16_16 (.ZN(mem_backbone_0_n_16_8), .A1(
      mem_backbone_0_ext_mem_din_sel[1]), .A2(pmem_dout[8]), .B1(
      mem_backbone_0_n_4), .B2(mem_backbone_0_per_dout_val[8]), .C1(
      mem_backbone_0_n_3), .C2(dmem_dout[8]));
  INV_X1_LVT mem_backbone_0_i_16_17 (.ZN(dbg_mem_din[8]), .A(
      mem_backbone_0_n_16_8));
  DFFR_X1_LVT \mem_backbone_0_per_dout_val_reg[7] (.Q(
      mem_backbone_0_per_dout_val[7]), .QN(), .CK(mclk), .D(per_dout_or[7]), .RN(
      mem_backbone_0_n_2));
  AOI222_X1_LVT mem_backbone_0_i_16_14 (.ZN(mem_backbone_0_n_16_7), .A1(
      mem_backbone_0_ext_mem_din_sel[1]), .A2(pmem_dout[7]), .B1(
      mem_backbone_0_n_4), .B2(mem_backbone_0_per_dout_val[7]), .C1(
      mem_backbone_0_n_3), .C2(dmem_dout[7]));
  INV_X1_LVT mem_backbone_0_i_16_15 (.ZN(dbg_mem_din[7]), .A(
      mem_backbone_0_n_16_7));
  DFFR_X1_LVT \mem_backbone_0_per_dout_val_reg[6] (.Q(
      mem_backbone_0_per_dout_val[6]), .QN(), .CK(mclk), .D(per_dout_or[6]), .RN(
      mem_backbone_0_n_2));
  AOI222_X1_LVT mem_backbone_0_i_16_12 (.ZN(mem_backbone_0_n_16_6), .A1(
      mem_backbone_0_ext_mem_din_sel[1]), .A2(pmem_dout[6]), .B1(
      mem_backbone_0_n_4), .B2(mem_backbone_0_per_dout_val[6]), .C1(
      mem_backbone_0_n_3), .C2(dmem_dout[6]));
  INV_X1_LVT mem_backbone_0_i_16_13 (.ZN(dbg_mem_din[6]), .A(
      mem_backbone_0_n_16_6));
  DFFR_X1_LVT \mem_backbone_0_per_dout_val_reg[5] (.Q(
      mem_backbone_0_per_dout_val[5]), .QN(), .CK(mclk), .D(per_dout_or[5]), .RN(
      mem_backbone_0_n_2));
  AOI222_X1_LVT mem_backbone_0_i_16_10 (.ZN(mem_backbone_0_n_16_5), .A1(
      mem_backbone_0_ext_mem_din_sel[1]), .A2(pmem_dout[5]), .B1(
      mem_backbone_0_n_4), .B2(mem_backbone_0_per_dout_val[5]), .C1(
      mem_backbone_0_n_3), .C2(dmem_dout[5]));
  INV_X1_LVT mem_backbone_0_i_16_11 (.ZN(dbg_mem_din[5]), .A(
      mem_backbone_0_n_16_5));
  DFFR_X1_LVT \mem_backbone_0_per_dout_val_reg[4] (.Q(
      mem_backbone_0_per_dout_val[4]), .QN(), .CK(mclk), .D(per_dout_or[4]), .RN(
      mem_backbone_0_n_2));
  AOI222_X1_LVT mem_backbone_0_i_16_8 (.ZN(mem_backbone_0_n_16_4), .A1(
      mem_backbone_0_ext_mem_din_sel[1]), .A2(pmem_dout[4]), .B1(
      mem_backbone_0_n_4), .B2(mem_backbone_0_per_dout_val[4]), .C1(
      mem_backbone_0_n_3), .C2(dmem_dout[4]));
  INV_X1_LVT mem_backbone_0_i_16_9 (.ZN(dbg_mem_din[4]), .A(
      mem_backbone_0_n_16_4));
  DFFR_X1_LVT \mem_backbone_0_per_dout_val_reg[3] (.Q(
      mem_backbone_0_per_dout_val[3]), .QN(), .CK(mclk), .D(per_dout_or[3]), .RN(
      mem_backbone_0_n_2));
  AOI222_X1_LVT mem_backbone_0_i_16_6 (.ZN(mem_backbone_0_n_16_3), .A1(
      mem_backbone_0_ext_mem_din_sel[1]), .A2(pmem_dout[3]), .B1(
      mem_backbone_0_n_4), .B2(mem_backbone_0_per_dout_val[3]), .C1(
      mem_backbone_0_n_3), .C2(dmem_dout[3]));
  INV_X1_LVT mem_backbone_0_i_16_7 (.ZN(dbg_mem_din[3]), .A(
      mem_backbone_0_n_16_3));
  DFFR_X1_LVT \mem_backbone_0_per_dout_val_reg[2] (.Q(
      mem_backbone_0_per_dout_val[2]), .QN(), .CK(mclk), .D(per_dout_or[2]), .RN(
      mem_backbone_0_n_2));
  AOI222_X1_LVT mem_backbone_0_i_16_4 (.ZN(mem_backbone_0_n_16_2), .A1(
      mem_backbone_0_ext_mem_din_sel[1]), .A2(pmem_dout[2]), .B1(
      mem_backbone_0_n_4), .B2(mem_backbone_0_per_dout_val[2]), .C1(
      mem_backbone_0_n_3), .C2(dmem_dout[2]));
  INV_X1_LVT mem_backbone_0_i_16_5 (.ZN(dbg_mem_din[2]), .A(
      mem_backbone_0_n_16_2));
  DFFR_X1_LVT \mem_backbone_0_per_dout_val_reg[1] (.Q(
      mem_backbone_0_per_dout_val[1]), .QN(), .CK(mclk), .D(per_dout_or[1]), .RN(
      mem_backbone_0_n_2));
  AOI222_X1_LVT mem_backbone_0_i_16_2 (.ZN(mem_backbone_0_n_16_1), .A1(
      mem_backbone_0_ext_mem_din_sel[1]), .A2(pmem_dout[1]), .B1(
      mem_backbone_0_n_4), .B2(mem_backbone_0_per_dout_val[1]), .C1(
      mem_backbone_0_n_3), .C2(dmem_dout[1]));
  INV_X1_LVT mem_backbone_0_i_16_3 (.ZN(dbg_mem_din[1]), .A(
      mem_backbone_0_n_16_1));
  DFFR_X1_LVT \mem_backbone_0_per_dout_val_reg[0] (.Q(
      mem_backbone_0_per_dout_val[0]), .QN(), .CK(mclk), .D(per_dout_or[0]), .RN(
      mem_backbone_0_n_2));
  AOI222_X1_LVT mem_backbone_0_i_16_0 (.ZN(mem_backbone_0_n_16_0), .A1(
      pmem_dout[0]), .A2(mem_backbone_0_ext_mem_din_sel[1]), .B1(
      mem_backbone_0_per_dout_val[0]), .B2(mem_backbone_0_n_4), .C1(dmem_dout[0]), 
      .C2(mem_backbone_0_n_3));
  INV_X1_LVT mem_backbone_0_i_16_1 (.ZN(dbg_mem_din[0]), .A(mem_backbone_0_n_16_0));
  INV_X1_LVT mem_backbone_0_i_19_0 (.ZN(mem_backbone_0_n_19_0), .A(
      mem_backbone_0_ext_mem_addr[11]));
  INV_X1_LVT mem_backbone_0_i_19_1 (.ZN(mem_backbone_0_n_19_1), .A(
      mem_backbone_0_ext_mem_addr[12]));
  INV_X1_LVT mem_backbone_0_i_19_2 (.ZN(mem_backbone_0_n_19_2), .A(
      mem_backbone_0_ext_mem_addr[13]));
  INV_X1_LVT mem_backbone_0_i_19_3 (.ZN(mem_backbone_0_n_19_3), .A(
      mem_backbone_0_ext_mem_addr[14]));
  NAND4_X1_LVT mem_backbone_0_i_19_4 (.ZN(mem_backbone_0_n_19_4), .A1(
      mem_backbone_0_n_19_0), .A2(mem_backbone_0_n_19_1), .A3(
      mem_backbone_0_n_19_2), .A4(mem_backbone_0_n_19_3));
  NOR4_X1_LVT mem_backbone_0_i_19_5 (.ZN(mem_backbone_0_n_19_5), .A1(
      mem_backbone_0_n_19_4), .A2(mem_backbone_0_ext_mem_addr[8]), .A3(
      mem_backbone_0_ext_mem_addr[9]), .A4(mem_backbone_0_ext_mem_addr[10]));
  AND2_X1_LVT mem_backbone_0_i_19_6 (.ZN(mem_backbone_0_n_19_6), .A1(
      mem_backbone_0_ext_mem_addr[8]), .A2(mem_backbone_0_ext_mem_addr[9]));
  NOR4_X1_LVT mem_backbone_0_i_19_7 (.ZN(mem_backbone_0_ext_dmem_sel), .A1(
      mem_backbone_0_n_19_4), .A2(mem_backbone_0_n_19_5), .A3(
      mem_backbone_0_n_19_6), .A4(mem_backbone_0_ext_mem_addr[10]));
  NAND2_X1_LVT mem_backbone_0_i_21_0 (.ZN(mem_backbone_0_n_21_0), .A1(
      mem_backbone_0_ext_mem_en), .A2(mem_backbone_0_ext_dmem_sel));
  OR4_X1_LVT mem_backbone_0_i_20_0 (.ZN(mem_backbone_0_n_20_0), .A1(eu_mab[12]), 
      .A2(eu_mab[13]), .A3(eu_mab[14]), .A4(eu_mab[15]));
  NOR4_X1_LVT mem_backbone_0_i_20_1 (.ZN(mem_backbone_0_n_20_1), .A1(
      mem_backbone_0_n_20_0), .A2(eu_mab[9]), .A3(eu_mab[10]), .A4(eu_mab[11]));
  AND2_X1_LVT mem_backbone_0_i_20_2 (.ZN(mem_backbone_0_n_20_2), .A1(eu_mab[9]), 
      .A2(eu_mab[10]));
  NOR4_X1_LVT mem_backbone_0_i_20_3 (.ZN(mem_backbone_0_n_20_3), .A1(
      mem_backbone_0_n_20_1), .A2(mem_backbone_0_n_20_2), .A3(eu_mab[11]), .A4(
      eu_mab[12]));
  INV_X1_LVT mem_backbone_0_i_20_4 (.ZN(mem_backbone_0_n_20_4), .A(eu_mb_en));
  NOR4_X1_LVT mem_backbone_0_i_20_5 (.ZN(mem_backbone_0_n_20_5), .A1(
      mem_backbone_0_n_20_4), .A2(eu_mab[13]), .A3(eu_mab[14]), .A4(eu_mab[15]));
  AND2_X1_LVT mem_backbone_0_i_20_6 (.ZN(mem_backbone_0_eu_dmem_en), .A1(
      mem_backbone_0_n_20_3), .A2(mem_backbone_0_n_20_5));
  NOR2_X1_LVT mem_backbone_0_i_21_1 (.ZN(mem_backbone_0_ext_dmem_en), .A1(
      mem_backbone_0_n_21_0), .A2(mem_backbone_0_eu_dmem_en));
  INV_X1_LVT mem_backbone_0_i_22_0 (.ZN(mem_backbone_0_n_22_0), .A(
      mem_backbone_0_ext_dmem_en));
  INV_X1_LVT mem_backbone_0_i_17_0 (.ZN(mem_backbone_0_n_5), .A(eu_mab[9]));
  INV_X1_LVT mem_backbone_0_i_18_0 (.ZN(mem_backbone_0_n_6), .A(
      mem_backbone_0_ext_mem_addr[8]));
  AOI22_X1_LVT mem_backbone_0_i_22_17 (.ZN(mem_backbone_0_n_22_9), .A1(
      mem_backbone_0_n_22_0), .A2(mem_backbone_0_n_5), .B1(
      mem_backbone_0_ext_dmem_en), .B2(mem_backbone_0_n_6));
  INV_X1_LVT mem_backbone_0_i_22_18 (.ZN(dmem_addr[8]), .A(mem_backbone_0_n_22_9));
  AOI22_X1_LVT mem_backbone_0_i_2_15 (.ZN(mem_backbone_0_n_2_8), .A1(
      mem_backbone_0_n_2_0), .A2(dma_addr[7]), .B1(dbg_mem_en), .B2(
      dbg_mem_addr[8]));
  INV_X1_LVT mem_backbone_0_i_2_16 (.ZN(mem_backbone_0_ext_mem_addr[7]), .A(
      mem_backbone_0_n_2_8));
  AOI22_X1_LVT mem_backbone_0_i_22_15 (.ZN(mem_backbone_0_n_22_8), .A1(
      mem_backbone_0_n_22_0), .A2(eu_mab[8]), .B1(mem_backbone_0_ext_dmem_en), 
      .B2(mem_backbone_0_ext_mem_addr[7]));
  INV_X1_LVT mem_backbone_0_i_22_16 (.ZN(dmem_addr[7]), .A(mem_backbone_0_n_22_8));
  AOI22_X1_LVT mem_backbone_0_i_2_13 (.ZN(mem_backbone_0_n_2_7), .A1(
      mem_backbone_0_n_2_0), .A2(dma_addr[6]), .B1(dbg_mem_en), .B2(
      dbg_mem_addr[7]));
  INV_X1_LVT mem_backbone_0_i_2_14 (.ZN(mem_backbone_0_ext_mem_addr[6]), .A(
      mem_backbone_0_n_2_7));
  AOI22_X1_LVT mem_backbone_0_i_22_13 (.ZN(mem_backbone_0_n_22_7), .A1(
      mem_backbone_0_n_22_0), .A2(eu_mab[7]), .B1(mem_backbone_0_ext_dmem_en), 
      .B2(mem_backbone_0_ext_mem_addr[6]));
  INV_X1_LVT mem_backbone_0_i_22_14 (.ZN(dmem_addr[6]), .A(mem_backbone_0_n_22_7));
  AOI22_X1_LVT mem_backbone_0_i_2_11 (.ZN(mem_backbone_0_n_2_6), .A1(
      mem_backbone_0_n_2_0), .A2(dma_addr[5]), .B1(dbg_mem_en), .B2(
      dbg_mem_addr[6]));
  INV_X1_LVT mem_backbone_0_i_2_12 (.ZN(mem_backbone_0_ext_mem_addr[5]), .A(
      mem_backbone_0_n_2_6));
  AOI22_X1_LVT mem_backbone_0_i_22_11 (.ZN(mem_backbone_0_n_22_6), .A1(
      mem_backbone_0_n_22_0), .A2(eu_mab[6]), .B1(mem_backbone_0_ext_dmem_en), 
      .B2(mem_backbone_0_ext_mem_addr[5]));
  INV_X1_LVT mem_backbone_0_i_22_12 (.ZN(dmem_addr[5]), .A(mem_backbone_0_n_22_6));
  AOI22_X1_LVT mem_backbone_0_i_2_9 (.ZN(mem_backbone_0_n_2_5), .A1(
      mem_backbone_0_n_2_0), .A2(dma_addr[4]), .B1(dbg_mem_en), .B2(
      dbg_mem_addr[5]));
  INV_X1_LVT mem_backbone_0_i_2_10 (.ZN(mem_backbone_0_ext_mem_addr[4]), .A(
      mem_backbone_0_n_2_5));
  AOI22_X1_LVT mem_backbone_0_i_22_9 (.ZN(mem_backbone_0_n_22_5), .A1(
      mem_backbone_0_n_22_0), .A2(eu_mab[5]), .B1(mem_backbone_0_ext_dmem_en), 
      .B2(mem_backbone_0_ext_mem_addr[4]));
  INV_X1_LVT mem_backbone_0_i_22_10 (.ZN(dmem_addr[4]), .A(mem_backbone_0_n_22_5));
  AOI22_X1_LVT mem_backbone_0_i_2_7 (.ZN(mem_backbone_0_n_2_4), .A1(
      mem_backbone_0_n_2_0), .A2(dma_addr[3]), .B1(dbg_mem_en), .B2(
      dbg_mem_addr[4]));
  INV_X1_LVT mem_backbone_0_i_2_8 (.ZN(mem_backbone_0_ext_mem_addr[3]), .A(
      mem_backbone_0_n_2_4));
  AOI22_X1_LVT mem_backbone_0_i_22_7 (.ZN(mem_backbone_0_n_22_4), .A1(
      mem_backbone_0_n_22_0), .A2(eu_mab[4]), .B1(mem_backbone_0_ext_dmem_en), 
      .B2(mem_backbone_0_ext_mem_addr[3]));
  INV_X1_LVT mem_backbone_0_i_22_8 (.ZN(dmem_addr[3]), .A(mem_backbone_0_n_22_4));
  AOI22_X1_LVT mem_backbone_0_i_2_5 (.ZN(mem_backbone_0_n_2_3), .A1(
      mem_backbone_0_n_2_0), .A2(dma_addr[2]), .B1(dbg_mem_en), .B2(
      dbg_mem_addr[3]));
  INV_X1_LVT mem_backbone_0_i_2_6 (.ZN(mem_backbone_0_ext_mem_addr[2]), .A(
      mem_backbone_0_n_2_3));
  AOI22_X1_LVT mem_backbone_0_i_22_5 (.ZN(mem_backbone_0_n_22_3), .A1(
      mem_backbone_0_n_22_0), .A2(eu_mab[3]), .B1(mem_backbone_0_ext_dmem_en), 
      .B2(mem_backbone_0_ext_mem_addr[2]));
  INV_X1_LVT mem_backbone_0_i_22_6 (.ZN(dmem_addr[2]), .A(mem_backbone_0_n_22_3));
  AOI22_X1_LVT mem_backbone_0_i_2_3 (.ZN(mem_backbone_0_n_2_2), .A1(
      mem_backbone_0_n_2_0), .A2(dma_addr[1]), .B1(dbg_mem_en), .B2(
      dbg_mem_addr[2]));
  INV_X1_LVT mem_backbone_0_i_2_4 (.ZN(mem_backbone_0_ext_mem_addr[1]), .A(
      mem_backbone_0_n_2_2));
  AOI22_X1_LVT mem_backbone_0_i_22_3 (.ZN(mem_backbone_0_n_22_2), .A1(
      mem_backbone_0_n_22_0), .A2(eu_mab[2]), .B1(mem_backbone_0_ext_dmem_en), 
      .B2(mem_backbone_0_ext_mem_addr[1]));
  INV_X1_LVT mem_backbone_0_i_22_4 (.ZN(dmem_addr[1]), .A(mem_backbone_0_n_22_2));
  AOI22_X1_LVT mem_backbone_0_i_2_1 (.ZN(mem_backbone_0_n_2_1), .A1(
      mem_backbone_0_n_2_0), .A2(dma_addr[0]), .B1(dbg_mem_addr[1]), .B2(
      dbg_mem_en));
  INV_X1_LVT mem_backbone_0_i_2_2 (.ZN(mem_backbone_0_ext_mem_addr[0]), .A(
      mem_backbone_0_n_2_1));
  AOI22_X1_LVT mem_backbone_0_i_22_1 (.ZN(mem_backbone_0_n_22_1), .A1(
      mem_backbone_0_n_22_0), .A2(eu_mab[1]), .B1(mem_backbone_0_ext_mem_addr[0]), 
      .B2(mem_backbone_0_ext_dmem_en));
  INV_X1_LVT mem_backbone_0_i_22_2 (.ZN(dmem_addr[0]), .A(mem_backbone_0_n_22_1));
  NOR2_X1_LVT mem_backbone_0_i_23_0 (.ZN(dmem_cen), .A1(
      mem_backbone_0_ext_dmem_en), .A2(mem_backbone_0_eu_dmem_en));
  INV_X1_LVT mem_backbone_0_i_25_0 (.ZN(mem_backbone_0_n_25_0), .A(
      mem_backbone_0_ext_dmem_en));
  INV_X1_LVT mem_backbone_0_i_24_0 (.ZN(mem_backbone_0_n_24_0), .A(dbg_mem_en));
  AOI22_X1_LVT mem_backbone_0_i_24_31 (.ZN(mem_backbone_0_n_24_16), .A1(
      mem_backbone_0_n_24_0), .A2(dma_din[15]), .B1(dbg_mem_en), .B2(
      dbg_mem_dout[15]));
  INV_X1_LVT mem_backbone_0_i_24_32 (.ZN(pmem_din[15]), .A(
      mem_backbone_0_n_24_16));
  AOI22_X1_LVT mem_backbone_0_i_25_31 (.ZN(mem_backbone_0_n_25_16), .A1(
      mem_backbone_0_n_25_0), .A2(eu_mdb_out[15]), .B1(
      mem_backbone_0_ext_dmem_en), .B2(pmem_din[15]));
  INV_X1_LVT mem_backbone_0_i_25_32 (.ZN(dmem_din[15]), .A(
      mem_backbone_0_n_25_16));
  AOI22_X1_LVT mem_backbone_0_i_24_29 (.ZN(mem_backbone_0_n_24_15), .A1(
      mem_backbone_0_n_24_0), .A2(dma_din[14]), .B1(dbg_mem_en), .B2(
      dbg_mem_dout[14]));
  INV_X1_LVT mem_backbone_0_i_24_30 (.ZN(pmem_din[14]), .A(
      mem_backbone_0_n_24_15));
  AOI22_X1_LVT mem_backbone_0_i_25_29 (.ZN(mem_backbone_0_n_25_15), .A1(
      mem_backbone_0_n_25_0), .A2(eu_mdb_out[14]), .B1(
      mem_backbone_0_ext_dmem_en), .B2(pmem_din[14]));
  INV_X1_LVT mem_backbone_0_i_25_30 (.ZN(dmem_din[14]), .A(
      mem_backbone_0_n_25_15));
  AOI22_X1_LVT mem_backbone_0_i_24_27 (.ZN(mem_backbone_0_n_24_14), .A1(
      mem_backbone_0_n_24_0), .A2(dma_din[13]), .B1(dbg_mem_en), .B2(
      dbg_mem_dout[13]));
  INV_X1_LVT mem_backbone_0_i_24_28 (.ZN(pmem_din[13]), .A(
      mem_backbone_0_n_24_14));
  AOI22_X1_LVT mem_backbone_0_i_25_27 (.ZN(mem_backbone_0_n_25_14), .A1(
      mem_backbone_0_n_25_0), .A2(eu_mdb_out[13]), .B1(
      mem_backbone_0_ext_dmem_en), .B2(pmem_din[13]));
  INV_X1_LVT mem_backbone_0_i_25_28 (.ZN(dmem_din[13]), .A(
      mem_backbone_0_n_25_14));
  AOI22_X1_LVT mem_backbone_0_i_24_25 (.ZN(mem_backbone_0_n_24_13), .A1(
      mem_backbone_0_n_24_0), .A2(dma_din[12]), .B1(dbg_mem_en), .B2(
      dbg_mem_dout[12]));
  INV_X1_LVT mem_backbone_0_i_24_26 (.ZN(pmem_din[12]), .A(
      mem_backbone_0_n_24_13));
  AOI22_X1_LVT mem_backbone_0_i_25_25 (.ZN(mem_backbone_0_n_25_13), .A1(
      mem_backbone_0_n_25_0), .A2(eu_mdb_out[12]), .B1(
      mem_backbone_0_ext_dmem_en), .B2(pmem_din[12]));
  INV_X1_LVT mem_backbone_0_i_25_26 (.ZN(dmem_din[12]), .A(
      mem_backbone_0_n_25_13));
  AOI22_X1_LVT mem_backbone_0_i_24_23 (.ZN(mem_backbone_0_n_24_12), .A1(
      mem_backbone_0_n_24_0), .A2(dma_din[11]), .B1(dbg_mem_en), .B2(
      dbg_mem_dout[11]));
  INV_X1_LVT mem_backbone_0_i_24_24 (.ZN(pmem_din[11]), .A(
      mem_backbone_0_n_24_12));
  AOI22_X1_LVT mem_backbone_0_i_25_23 (.ZN(mem_backbone_0_n_25_12), .A1(
      mem_backbone_0_n_25_0), .A2(eu_mdb_out[11]), .B1(
      mem_backbone_0_ext_dmem_en), .B2(pmem_din[11]));
  INV_X1_LVT mem_backbone_0_i_25_24 (.ZN(dmem_din[11]), .A(
      mem_backbone_0_n_25_12));
  AOI22_X1_LVT mem_backbone_0_i_24_21 (.ZN(mem_backbone_0_n_24_11), .A1(
      mem_backbone_0_n_24_0), .A2(dma_din[10]), .B1(dbg_mem_en), .B2(
      dbg_mem_dout[10]));
  INV_X1_LVT mem_backbone_0_i_24_22 (.ZN(pmem_din[10]), .A(
      mem_backbone_0_n_24_11));
  AOI22_X1_LVT mem_backbone_0_i_25_21 (.ZN(mem_backbone_0_n_25_11), .A1(
      mem_backbone_0_n_25_0), .A2(eu_mdb_out[10]), .B1(
      mem_backbone_0_ext_dmem_en), .B2(pmem_din[10]));
  INV_X1_LVT mem_backbone_0_i_25_22 (.ZN(dmem_din[10]), .A(
      mem_backbone_0_n_25_11));
  AOI22_X1_LVT mem_backbone_0_i_24_19 (.ZN(mem_backbone_0_n_24_10), .A1(
      mem_backbone_0_n_24_0), .A2(dma_din[9]), .B1(dbg_mem_en), .B2(
      dbg_mem_dout[9]));
  INV_X1_LVT mem_backbone_0_i_24_20 (.ZN(pmem_din[9]), .A(mem_backbone_0_n_24_10));
  AOI22_X1_LVT mem_backbone_0_i_25_19 (.ZN(mem_backbone_0_n_25_10), .A1(
      mem_backbone_0_n_25_0), .A2(eu_mdb_out[9]), .B1(mem_backbone_0_ext_dmem_en), 
      .B2(pmem_din[9]));
  INV_X1_LVT mem_backbone_0_i_25_20 (.ZN(dmem_din[9]), .A(mem_backbone_0_n_25_10));
  AOI22_X1_LVT mem_backbone_0_i_24_17 (.ZN(mem_backbone_0_n_24_9), .A1(
      mem_backbone_0_n_24_0), .A2(dma_din[8]), .B1(dbg_mem_en), .B2(
      dbg_mem_dout[8]));
  INV_X1_LVT mem_backbone_0_i_24_18 (.ZN(pmem_din[8]), .A(mem_backbone_0_n_24_9));
  AOI22_X1_LVT mem_backbone_0_i_25_17 (.ZN(mem_backbone_0_n_25_9), .A1(
      mem_backbone_0_n_25_0), .A2(eu_mdb_out[8]), .B1(mem_backbone_0_ext_dmem_en), 
      .B2(pmem_din[8]));
  INV_X1_LVT mem_backbone_0_i_25_18 (.ZN(dmem_din[8]), .A(mem_backbone_0_n_25_9));
  AOI22_X1_LVT mem_backbone_0_i_24_15 (.ZN(mem_backbone_0_n_24_8), .A1(
      mem_backbone_0_n_24_0), .A2(dma_din[7]), .B1(dbg_mem_en), .B2(
      dbg_mem_dout[7]));
  INV_X1_LVT mem_backbone_0_i_24_16 (.ZN(pmem_din[7]), .A(mem_backbone_0_n_24_8));
  AOI22_X1_LVT mem_backbone_0_i_25_15 (.ZN(mem_backbone_0_n_25_8), .A1(
      mem_backbone_0_n_25_0), .A2(eu_mdb_out[7]), .B1(mem_backbone_0_ext_dmem_en), 
      .B2(pmem_din[7]));
  INV_X1_LVT mem_backbone_0_i_25_16 (.ZN(dmem_din[7]), .A(mem_backbone_0_n_25_8));
  AOI22_X1_LVT mem_backbone_0_i_24_13 (.ZN(mem_backbone_0_n_24_7), .A1(
      mem_backbone_0_n_24_0), .A2(dma_din[6]), .B1(dbg_mem_en), .B2(
      dbg_mem_dout[6]));
  INV_X1_LVT mem_backbone_0_i_24_14 (.ZN(pmem_din[6]), .A(mem_backbone_0_n_24_7));
  AOI22_X1_LVT mem_backbone_0_i_25_13 (.ZN(mem_backbone_0_n_25_7), .A1(
      mem_backbone_0_n_25_0), .A2(eu_mdb_out[6]), .B1(mem_backbone_0_ext_dmem_en), 
      .B2(pmem_din[6]));
  INV_X1_LVT mem_backbone_0_i_25_14 (.ZN(dmem_din[6]), .A(mem_backbone_0_n_25_7));
  AOI22_X1_LVT mem_backbone_0_i_24_11 (.ZN(mem_backbone_0_n_24_6), .A1(
      mem_backbone_0_n_24_0), .A2(dma_din[5]), .B1(dbg_mem_en), .B2(
      dbg_mem_dout[5]));
  INV_X1_LVT mem_backbone_0_i_24_12 (.ZN(pmem_din[5]), .A(mem_backbone_0_n_24_6));
  AOI22_X1_LVT mem_backbone_0_i_25_11 (.ZN(mem_backbone_0_n_25_6), .A1(
      mem_backbone_0_n_25_0), .A2(eu_mdb_out[5]), .B1(mem_backbone_0_ext_dmem_en), 
      .B2(pmem_din[5]));
  INV_X1_LVT mem_backbone_0_i_25_12 (.ZN(dmem_din[5]), .A(mem_backbone_0_n_25_6));
  AOI22_X1_LVT mem_backbone_0_i_24_9 (.ZN(mem_backbone_0_n_24_5), .A1(
      mem_backbone_0_n_24_0), .A2(dma_din[4]), .B1(dbg_mem_en), .B2(
      dbg_mem_dout[4]));
  INV_X1_LVT mem_backbone_0_i_24_10 (.ZN(pmem_din[4]), .A(mem_backbone_0_n_24_5));
  AOI22_X1_LVT mem_backbone_0_i_25_9 (.ZN(mem_backbone_0_n_25_5), .A1(
      mem_backbone_0_n_25_0), .A2(eu_mdb_out[4]), .B1(mem_backbone_0_ext_dmem_en), 
      .B2(pmem_din[4]));
  INV_X1_LVT mem_backbone_0_i_25_10 (.ZN(dmem_din[4]), .A(mem_backbone_0_n_25_5));
  AOI22_X1_LVT mem_backbone_0_i_24_7 (.ZN(mem_backbone_0_n_24_4), .A1(
      mem_backbone_0_n_24_0), .A2(dma_din[3]), .B1(dbg_mem_en), .B2(
      dbg_mem_dout[3]));
  INV_X1_LVT mem_backbone_0_i_24_8 (.ZN(pmem_din[3]), .A(mem_backbone_0_n_24_4));
  AOI22_X1_LVT mem_backbone_0_i_25_7 (.ZN(mem_backbone_0_n_25_4), .A1(
      mem_backbone_0_n_25_0), .A2(eu_mdb_out[3]), .B1(mem_backbone_0_ext_dmem_en), 
      .B2(pmem_din[3]));
  INV_X1_LVT mem_backbone_0_i_25_8 (.ZN(dmem_din[3]), .A(mem_backbone_0_n_25_4));
  AOI22_X1_LVT mem_backbone_0_i_24_5 (.ZN(mem_backbone_0_n_24_3), .A1(
      mem_backbone_0_n_24_0), .A2(dma_din[2]), .B1(dbg_mem_en), .B2(
      dbg_mem_dout[2]));
  INV_X1_LVT mem_backbone_0_i_24_6 (.ZN(pmem_din[2]), .A(mem_backbone_0_n_24_3));
  AOI22_X1_LVT mem_backbone_0_i_25_5 (.ZN(mem_backbone_0_n_25_3), .A1(
      mem_backbone_0_n_25_0), .A2(eu_mdb_out[2]), .B1(mem_backbone_0_ext_dmem_en), 
      .B2(pmem_din[2]));
  INV_X1_LVT mem_backbone_0_i_25_6 (.ZN(dmem_din[2]), .A(mem_backbone_0_n_25_3));
  AOI22_X1_LVT mem_backbone_0_i_24_3 (.ZN(mem_backbone_0_n_24_2), .A1(
      mem_backbone_0_n_24_0), .A2(dma_din[1]), .B1(dbg_mem_en), .B2(
      dbg_mem_dout[1]));
  INV_X1_LVT mem_backbone_0_i_24_4 (.ZN(pmem_din[1]), .A(mem_backbone_0_n_24_2));
  AOI22_X1_LVT mem_backbone_0_i_25_3 (.ZN(mem_backbone_0_n_25_2), .A1(
      mem_backbone_0_n_25_0), .A2(eu_mdb_out[1]), .B1(mem_backbone_0_ext_dmem_en), 
      .B2(pmem_din[1]));
  INV_X1_LVT mem_backbone_0_i_25_4 (.ZN(dmem_din[1]), .A(mem_backbone_0_n_25_2));
  AOI22_X1_LVT mem_backbone_0_i_24_1 (.ZN(mem_backbone_0_n_24_1), .A1(
      mem_backbone_0_n_24_0), .A2(dma_din[0]), .B1(dbg_mem_dout[0]), .B2(
      dbg_mem_en));
  INV_X1_LVT mem_backbone_0_i_24_2 (.ZN(pmem_din[0]), .A(mem_backbone_0_n_24_1));
  AOI22_X1_LVT mem_backbone_0_i_25_1 (.ZN(mem_backbone_0_n_25_1), .A1(
      mem_backbone_0_n_25_0), .A2(eu_mdb_out[0]), .B1(pmem_din[0]), .B2(
      mem_backbone_0_ext_dmem_en));
  INV_X1_LVT mem_backbone_0_i_25_2 (.ZN(dmem_din[0]), .A(mem_backbone_0_n_25_1));
  INV_X1_LVT mem_backbone_0_i_29_0 (.ZN(mem_backbone_0_n_29_0), .A(
      mem_backbone_0_ext_dmem_en));
  INV_X1_LVT mem_backbone_0_i_26_1 (.ZN(mem_backbone_0_n_8), .A(eu_mb_wr[1]));
  INV_X1_LVT mem_backbone_0_i_27_0 (.ZN(mem_backbone_0_n_27_0), .A(dbg_mem_en));
  AOI22_X1_LVT mem_backbone_0_i_27_3 (.ZN(mem_backbone_0_n_27_2), .A1(
      mem_backbone_0_n_27_0), .A2(dma_we[1]), .B1(dbg_mem_en), .B2(dbg_mem_wr[1]));
  INV_X1_LVT mem_backbone_0_i_27_4 (.ZN(mem_backbone_0_ext_mem_wr[1]), .A(
      mem_backbone_0_n_27_2));
  INV_X1_LVT mem_backbone_0_i_28_1 (.ZN(mem_backbone_0_n_10), .A(
      mem_backbone_0_ext_mem_wr[1]));
  AOI22_X1_LVT mem_backbone_0_i_29_3 (.ZN(mem_backbone_0_n_29_2), .A1(
      mem_backbone_0_n_29_0), .A2(mem_backbone_0_n_8), .B1(
      mem_backbone_0_ext_dmem_en), .B2(mem_backbone_0_n_10));
  INV_X1_LVT mem_backbone_0_i_29_4 (.ZN(dmem_wen[1]), .A(mem_backbone_0_n_29_2));
  INV_X1_LVT mem_backbone_0_i_26_0 (.ZN(mem_backbone_0_n_7), .A(eu_mb_wr[0]));
  AOI22_X1_LVT mem_backbone_0_i_27_1 (.ZN(mem_backbone_0_n_27_1), .A1(
      mem_backbone_0_n_27_0), .A2(dma_we[0]), .B1(dbg_mem_wr[0]), .B2(dbg_mem_en));
  INV_X1_LVT mem_backbone_0_i_27_2 (.ZN(mem_backbone_0_ext_mem_wr[0]), .A(
      mem_backbone_0_n_27_1));
  INV_X1_LVT mem_backbone_0_i_28_0 (.ZN(mem_backbone_0_n_9), .A(
      mem_backbone_0_ext_mem_wr[0]));
  AOI22_X1_LVT mem_backbone_0_i_29_1 (.ZN(mem_backbone_0_n_29_1), .A1(
      mem_backbone_0_n_29_0), .A2(mem_backbone_0_n_7), .B1(mem_backbone_0_n_9), 
      .B2(mem_backbone_0_ext_dmem_en));
  INV_X1_LVT mem_backbone_0_i_29_2 (.ZN(dmem_wen[0]), .A(mem_backbone_0_n_29_1));
  DFFR_X1_LVT \mem_backbone_0_eu_mdb_in_sel_reg[1] (.Q(
      mem_backbone_0_eu_mdb_in_sel[1]), .QN(), .CK(mclk), .D(
      mem_backbone_0_eu_pmem_en), .RN(mem_backbone_0_n_2));
  DFFR_X1_LVT \mem_backbone_0_eu_mdb_in_sel_reg[0] (.Q(
      mem_backbone_0_eu_mdb_in_sel[0]), .QN(), .CK(mclk), .D(
      mem_backbone_0_eu_per_en), .RN(mem_backbone_0_n_2));
  INV_X1_LVT mem_backbone_0_i_31_1 (.ZN(mem_backbone_0_n_31_0), .A(
      mem_backbone_0_eu_mdb_in_sel[0]));
  NOR2_X1_LVT mem_backbone_0_i_31_2 (.ZN(mem_backbone_0_n_12), .A1(
      mem_backbone_0_n_31_0), .A2(mem_backbone_0_eu_mdb_in_sel[1]));
  NOR2_X1_LVT mem_backbone_0_i_31_0 (.ZN(mem_backbone_0_n_11), .A1(
      mem_backbone_0_eu_mdb_in_sel[0]), .A2(mem_backbone_0_eu_mdb_in_sel[1]));
  AOI222_X1_LVT mem_backbone_0_i_32_30 (.ZN(mem_backbone_0_n_32_15), .A1(
      mem_backbone_0_eu_mdb_in_sel[1]), .A2(pmem_dout[15]), .B1(
      mem_backbone_0_n_12), .B2(mem_backbone_0_per_dout_val[15]), .C1(
      mem_backbone_0_n_11), .C2(dmem_dout[15]));
  INV_X1_LVT mem_backbone_0_i_32_31 (.ZN(eu_mdb_in[15]), .A(
      mem_backbone_0_n_32_15));
  AOI222_X1_LVT mem_backbone_0_i_32_28 (.ZN(mem_backbone_0_n_32_14), .A1(
      mem_backbone_0_eu_mdb_in_sel[1]), .A2(pmem_dout[14]), .B1(
      mem_backbone_0_n_12), .B2(mem_backbone_0_per_dout_val[14]), .C1(
      mem_backbone_0_n_11), .C2(dmem_dout[14]));
  INV_X1_LVT mem_backbone_0_i_32_29 (.ZN(eu_mdb_in[14]), .A(
      mem_backbone_0_n_32_14));
  AOI222_X1_LVT mem_backbone_0_i_32_26 (.ZN(mem_backbone_0_n_32_13), .A1(
      mem_backbone_0_eu_mdb_in_sel[1]), .A2(pmem_dout[13]), .B1(
      mem_backbone_0_n_12), .B2(mem_backbone_0_per_dout_val[13]), .C1(
      mem_backbone_0_n_11), .C2(dmem_dout[13]));
  INV_X1_LVT mem_backbone_0_i_32_27 (.ZN(eu_mdb_in[13]), .A(
      mem_backbone_0_n_32_13));
  AOI222_X1_LVT mem_backbone_0_i_32_24 (.ZN(mem_backbone_0_n_32_12), .A1(
      mem_backbone_0_eu_mdb_in_sel[1]), .A2(pmem_dout[12]), .B1(
      mem_backbone_0_n_12), .B2(mem_backbone_0_per_dout_val[12]), .C1(
      mem_backbone_0_n_11), .C2(dmem_dout[12]));
  INV_X1_LVT mem_backbone_0_i_32_25 (.ZN(eu_mdb_in[12]), .A(
      mem_backbone_0_n_32_12));
  AOI222_X1_LVT mem_backbone_0_i_32_22 (.ZN(mem_backbone_0_n_32_11), .A1(
      mem_backbone_0_eu_mdb_in_sel[1]), .A2(pmem_dout[11]), .B1(
      mem_backbone_0_n_12), .B2(mem_backbone_0_per_dout_val[11]), .C1(
      mem_backbone_0_n_11), .C2(dmem_dout[11]));
  INV_X1_LVT mem_backbone_0_i_32_23 (.ZN(eu_mdb_in[11]), .A(
      mem_backbone_0_n_32_11));
  AOI222_X1_LVT mem_backbone_0_i_32_20 (.ZN(mem_backbone_0_n_32_10), .A1(
      mem_backbone_0_eu_mdb_in_sel[1]), .A2(pmem_dout[10]), .B1(
      mem_backbone_0_n_12), .B2(mem_backbone_0_per_dout_val[10]), .C1(
      mem_backbone_0_n_11), .C2(dmem_dout[10]));
  INV_X1_LVT mem_backbone_0_i_32_21 (.ZN(eu_mdb_in[10]), .A(
      mem_backbone_0_n_32_10));
  AOI222_X1_LVT mem_backbone_0_i_32_18 (.ZN(mem_backbone_0_n_32_9), .A1(
      mem_backbone_0_eu_mdb_in_sel[1]), .A2(pmem_dout[9]), .B1(
      mem_backbone_0_n_12), .B2(mem_backbone_0_per_dout_val[9]), .C1(
      mem_backbone_0_n_11), .C2(dmem_dout[9]));
  INV_X1_LVT mem_backbone_0_i_32_19 (.ZN(eu_mdb_in[9]), .A(mem_backbone_0_n_32_9));
  AOI222_X1_LVT mem_backbone_0_i_32_16 (.ZN(mem_backbone_0_n_32_8), .A1(
      mem_backbone_0_eu_mdb_in_sel[1]), .A2(pmem_dout[8]), .B1(
      mem_backbone_0_n_12), .B2(mem_backbone_0_per_dout_val[8]), .C1(
      mem_backbone_0_n_11), .C2(dmem_dout[8]));
  INV_X1_LVT mem_backbone_0_i_32_17 (.ZN(eu_mdb_in[8]), .A(mem_backbone_0_n_32_8));
  AOI222_X1_LVT mem_backbone_0_i_32_14 (.ZN(mem_backbone_0_n_32_7), .A1(
      mem_backbone_0_eu_mdb_in_sel[1]), .A2(pmem_dout[7]), .B1(
      mem_backbone_0_n_12), .B2(mem_backbone_0_per_dout_val[7]), .C1(
      mem_backbone_0_n_11), .C2(dmem_dout[7]));
  INV_X1_LVT mem_backbone_0_i_32_15 (.ZN(eu_mdb_in[7]), .A(mem_backbone_0_n_32_7));
  AOI222_X1_LVT mem_backbone_0_i_32_12 (.ZN(mem_backbone_0_n_32_6), .A1(
      mem_backbone_0_eu_mdb_in_sel[1]), .A2(pmem_dout[6]), .B1(
      mem_backbone_0_n_12), .B2(mem_backbone_0_per_dout_val[6]), .C1(
      mem_backbone_0_n_11), .C2(dmem_dout[6]));
  INV_X1_LVT mem_backbone_0_i_32_13 (.ZN(eu_mdb_in[6]), .A(mem_backbone_0_n_32_6));
  AOI222_X1_LVT mem_backbone_0_i_32_10 (.ZN(mem_backbone_0_n_32_5), .A1(
      mem_backbone_0_eu_mdb_in_sel[1]), .A2(pmem_dout[5]), .B1(
      mem_backbone_0_n_12), .B2(mem_backbone_0_per_dout_val[5]), .C1(
      mem_backbone_0_n_11), .C2(dmem_dout[5]));
  INV_X1_LVT mem_backbone_0_i_32_11 (.ZN(eu_mdb_in[5]), .A(mem_backbone_0_n_32_5));
  AOI222_X1_LVT mem_backbone_0_i_32_8 (.ZN(mem_backbone_0_n_32_4), .A1(
      mem_backbone_0_eu_mdb_in_sel[1]), .A2(pmem_dout[4]), .B1(
      mem_backbone_0_n_12), .B2(mem_backbone_0_per_dout_val[4]), .C1(
      mem_backbone_0_n_11), .C2(dmem_dout[4]));
  INV_X1_LVT mem_backbone_0_i_32_9 (.ZN(eu_mdb_in[4]), .A(mem_backbone_0_n_32_4));
  AOI222_X1_LVT mem_backbone_0_i_32_6 (.ZN(mem_backbone_0_n_32_3), .A1(
      mem_backbone_0_eu_mdb_in_sel[1]), .A2(pmem_dout[3]), .B1(
      mem_backbone_0_n_12), .B2(mem_backbone_0_per_dout_val[3]), .C1(
      mem_backbone_0_n_11), .C2(dmem_dout[3]));
  INV_X1_LVT mem_backbone_0_i_32_7 (.ZN(eu_mdb_in[3]), .A(mem_backbone_0_n_32_3));
  AOI222_X1_LVT mem_backbone_0_i_32_4 (.ZN(mem_backbone_0_n_32_2), .A1(
      mem_backbone_0_eu_mdb_in_sel[1]), .A2(pmem_dout[2]), .B1(
      mem_backbone_0_n_12), .B2(mem_backbone_0_per_dout_val[2]), .C1(
      mem_backbone_0_n_11), .C2(dmem_dout[2]));
  INV_X1_LVT mem_backbone_0_i_32_5 (.ZN(eu_mdb_in[2]), .A(mem_backbone_0_n_32_2));
  AOI222_X1_LVT mem_backbone_0_i_32_2 (.ZN(mem_backbone_0_n_32_1), .A1(
      mem_backbone_0_eu_mdb_in_sel[1]), .A2(pmem_dout[1]), .B1(
      mem_backbone_0_n_12), .B2(mem_backbone_0_per_dout_val[1]), .C1(
      mem_backbone_0_n_11), .C2(dmem_dout[1]));
  INV_X1_LVT mem_backbone_0_i_32_3 (.ZN(eu_mdb_in[1]), .A(mem_backbone_0_n_32_1));
  AOI222_X1_LVT mem_backbone_0_i_32_0 (.ZN(mem_backbone_0_n_32_0), .A1(
      pmem_dout[0]), .A2(mem_backbone_0_eu_mdb_in_sel[1]), .B1(
      mem_backbone_0_per_dout_val[0]), .B2(mem_backbone_0_n_12), .C1(dmem_dout[0]), 
      .C2(mem_backbone_0_n_11));
  INV_X1_LVT mem_backbone_0_i_32_1 (.ZN(eu_mdb_in[0]), .A(mem_backbone_0_n_32_0));
  DFFR_X1_LVT mem_backbone_0_fe_pmem_en_dly_reg (.Q(
      mem_backbone_0_fe_pmem_en_dly), .QN(), .CK(mclk), .D(
      mem_backbone_0_fe_pmem_en), .RN(mem_backbone_0_n_2));
  NAND2_X1_LVT mem_backbone_0_i_33_0 (.ZN(mem_backbone_0_n_33_0), .A1(
      mem_backbone_0_n_0), .A2(mem_backbone_0_fe_pmem_en_dly));
  NOR2_X1_LVT mem_backbone_0_i_33_1 (.ZN(mem_backbone_0_fe_pmem_save), .A1(
      mem_backbone_0_n_33_0), .A2(cpu_halt_st));
  INV_X1_LVT mem_backbone_0_i_35_0 (.ZN(mem_backbone_0_n_35_0), .A(cpu_halt_st));
  INV_X1_LVT mem_backbone_0_i_35_1 (.ZN(mem_backbone_0_n_35_1), .A(
      mem_backbone_0_fe_pmem_en));
  OAI21_X1_LVT mem_backbone_0_i_35_2 (.ZN(mem_backbone_0_fe_pmem_restore), .A(
      mem_backbone_0_n_35_0), .B1(mem_backbone_0_n_35_1), .B2(
      mem_backbone_0_fe_pmem_en_dly));
  INV_X1_LVT mem_backbone_0_i_37_1 (.ZN(mem_backbone_0_n_37_1), .A(
      mem_backbone_0_fe_pmem_restore));
  INV_X1_LVT mem_backbone_0_i_37_0 (.ZN(mem_backbone_0_n_37_0), .A(
      mem_backbone_0_fe_pmem_save));
  NAND2_X1_LVT mem_backbone_0_i_37_2 (.ZN(mem_backbone_0_n_15), .A1(
      mem_backbone_0_n_37_1), .A2(mem_backbone_0_n_37_0));
  CLKGATETST_X1_LVT mem_backbone_0_clk_gate_pmem_dout_bckup_sel_reg (.GCK(
      mem_backbone_0_n_14), .CK(mclk), .E(mem_backbone_0_n_15), .SE(1'b0));
  DFFR_X1_LVT mem_backbone_0_pmem_dout_bckup_sel_reg (.Q(
      mem_backbone_0_pmem_dout_bckup_sel), .QN(), .CK(mem_backbone_0_n_14), .D(
      mem_backbone_0_fe_pmem_save), .RN(mem_backbone_0_n_2));
  INV_X1_LVT mem_backbone_0_i_39_0 (.ZN(mem_backbone_0_n_39_0), .A(
      mem_backbone_0_pmem_dout_bckup_sel));
  CLKGATETST_X1_LVT mem_backbone_0_clk_gate_pmem_dout_bckup_reg (.GCK(
      mem_backbone_0_n_13), .CK(mclk), .E(mem_backbone_0_fe_pmem_save), .SE(1'b0));
  DFFR_X1_LVT \mem_backbone_0_pmem_dout_bckup_reg[15] (.Q(
      mem_backbone_0_pmem_dout_bckup[15]), .QN(), .CK(mem_backbone_0_n_13), .D(
      pmem_dout[15]), .RN(mem_backbone_0_n_2));
  AOI22_X1_LVT mem_backbone_0_i_39_31 (.ZN(mem_backbone_0_n_39_16), .A1(
      mem_backbone_0_n_39_0), .A2(pmem_dout[15]), .B1(
      mem_backbone_0_pmem_dout_bckup_sel), .B2(
      mem_backbone_0_pmem_dout_bckup[15]));
  INV_X1_LVT mem_backbone_0_i_39_32 (.ZN(fe_mdb_in[15]), .A(
      mem_backbone_0_n_39_16));
  DFFR_X1_LVT \mem_backbone_0_pmem_dout_bckup_reg[14] (.Q(
      mem_backbone_0_pmem_dout_bckup[14]), .QN(), .CK(mem_backbone_0_n_13), .D(
      pmem_dout[14]), .RN(mem_backbone_0_n_2));
  AOI22_X1_LVT mem_backbone_0_i_39_29 (.ZN(mem_backbone_0_n_39_15), .A1(
      mem_backbone_0_n_39_0), .A2(pmem_dout[14]), .B1(
      mem_backbone_0_pmem_dout_bckup_sel), .B2(
      mem_backbone_0_pmem_dout_bckup[14]));
  INV_X1_LVT mem_backbone_0_i_39_30 (.ZN(fe_mdb_in[14]), .A(
      mem_backbone_0_n_39_15));
  DFFR_X1_LVT \mem_backbone_0_pmem_dout_bckup_reg[13] (.Q(
      mem_backbone_0_pmem_dout_bckup[13]), .QN(), .CK(mem_backbone_0_n_13), .D(
      pmem_dout[13]), .RN(mem_backbone_0_n_2));
  AOI22_X1_LVT mem_backbone_0_i_39_27 (.ZN(mem_backbone_0_n_39_14), .A1(
      mem_backbone_0_n_39_0), .A2(pmem_dout[13]), .B1(
      mem_backbone_0_pmem_dout_bckup_sel), .B2(
      mem_backbone_0_pmem_dout_bckup[13]));
  INV_X1_LVT mem_backbone_0_i_39_28 (.ZN(fe_mdb_in[13]), .A(
      mem_backbone_0_n_39_14));
  DFFR_X1_LVT \mem_backbone_0_pmem_dout_bckup_reg[12] (.Q(
      mem_backbone_0_pmem_dout_bckup[12]), .QN(), .CK(mem_backbone_0_n_13), .D(
      pmem_dout[12]), .RN(mem_backbone_0_n_2));
  AOI22_X1_LVT mem_backbone_0_i_39_25 (.ZN(mem_backbone_0_n_39_13), .A1(
      mem_backbone_0_n_39_0), .A2(pmem_dout[12]), .B1(
      mem_backbone_0_pmem_dout_bckup_sel), .B2(
      mem_backbone_0_pmem_dout_bckup[12]));
  INV_X1_LVT mem_backbone_0_i_39_26 (.ZN(fe_mdb_in[12]), .A(
      mem_backbone_0_n_39_13));
  DFFR_X1_LVT \mem_backbone_0_pmem_dout_bckup_reg[11] (.Q(
      mem_backbone_0_pmem_dout_bckup[11]), .QN(), .CK(mem_backbone_0_n_13), .D(
      pmem_dout[11]), .RN(mem_backbone_0_n_2));
  AOI22_X1_LVT mem_backbone_0_i_39_23 (.ZN(mem_backbone_0_n_39_12), .A1(
      mem_backbone_0_n_39_0), .A2(pmem_dout[11]), .B1(
      mem_backbone_0_pmem_dout_bckup_sel), .B2(
      mem_backbone_0_pmem_dout_bckup[11]));
  INV_X1_LVT mem_backbone_0_i_39_24 (.ZN(fe_mdb_in[11]), .A(
      mem_backbone_0_n_39_12));
  DFFR_X1_LVT \mem_backbone_0_pmem_dout_bckup_reg[10] (.Q(
      mem_backbone_0_pmem_dout_bckup[10]), .QN(), .CK(mem_backbone_0_n_13), .D(
      pmem_dout[10]), .RN(mem_backbone_0_n_2));
  AOI22_X1_LVT mem_backbone_0_i_39_21 (.ZN(mem_backbone_0_n_39_11), .A1(
      mem_backbone_0_n_39_0), .A2(pmem_dout[10]), .B1(
      mem_backbone_0_pmem_dout_bckup_sel), .B2(
      mem_backbone_0_pmem_dout_bckup[10]));
  INV_X1_LVT mem_backbone_0_i_39_22 (.ZN(fe_mdb_in[10]), .A(
      mem_backbone_0_n_39_11));
  DFFR_X1_LVT \mem_backbone_0_pmem_dout_bckup_reg[9] (.Q(
      mem_backbone_0_pmem_dout_bckup[9]), .QN(), .CK(mem_backbone_0_n_13), .D(
      pmem_dout[9]), .RN(mem_backbone_0_n_2));
  AOI22_X1_LVT mem_backbone_0_i_39_19 (.ZN(mem_backbone_0_n_39_10), .A1(
      mem_backbone_0_n_39_0), .A2(pmem_dout[9]), .B1(
      mem_backbone_0_pmem_dout_bckup_sel), .B2(mem_backbone_0_pmem_dout_bckup[9]));
  INV_X1_LVT mem_backbone_0_i_39_20 (.ZN(fe_mdb_in[9]), .A(
      mem_backbone_0_n_39_10));
  DFFR_X1_LVT \mem_backbone_0_pmem_dout_bckup_reg[8] (.Q(
      mem_backbone_0_pmem_dout_bckup[8]), .QN(), .CK(mem_backbone_0_n_13), .D(
      pmem_dout[8]), .RN(mem_backbone_0_n_2));
  AOI22_X1_LVT mem_backbone_0_i_39_17 (.ZN(mem_backbone_0_n_39_9), .A1(
      mem_backbone_0_n_39_0), .A2(pmem_dout[8]), .B1(
      mem_backbone_0_pmem_dout_bckup_sel), .B2(mem_backbone_0_pmem_dout_bckup[8]));
  INV_X1_LVT mem_backbone_0_i_39_18 (.ZN(fe_mdb_in[8]), .A(mem_backbone_0_n_39_9));
  DFFR_X1_LVT \mem_backbone_0_pmem_dout_bckup_reg[7] (.Q(
      mem_backbone_0_pmem_dout_bckup[7]), .QN(), .CK(mem_backbone_0_n_13), .D(
      pmem_dout[7]), .RN(mem_backbone_0_n_2));
  AOI22_X1_LVT mem_backbone_0_i_39_15 (.ZN(mem_backbone_0_n_39_8), .A1(
      mem_backbone_0_n_39_0), .A2(pmem_dout[7]), .B1(
      mem_backbone_0_pmem_dout_bckup_sel), .B2(mem_backbone_0_pmem_dout_bckup[7]));
  INV_X1_LVT mem_backbone_0_i_39_16 (.ZN(fe_mdb_in[7]), .A(mem_backbone_0_n_39_8));
  DFFR_X1_LVT \mem_backbone_0_pmem_dout_bckup_reg[6] (.Q(
      mem_backbone_0_pmem_dout_bckup[6]), .QN(), .CK(mem_backbone_0_n_13), .D(
      pmem_dout[6]), .RN(mem_backbone_0_n_2));
  AOI22_X1_LVT mem_backbone_0_i_39_13 (.ZN(mem_backbone_0_n_39_7), .A1(
      mem_backbone_0_n_39_0), .A2(pmem_dout[6]), .B1(
      mem_backbone_0_pmem_dout_bckup_sel), .B2(mem_backbone_0_pmem_dout_bckup[6]));
  INV_X1_LVT mem_backbone_0_i_39_14 (.ZN(fe_mdb_in[6]), .A(mem_backbone_0_n_39_7));
  DFFR_X1_LVT \mem_backbone_0_pmem_dout_bckup_reg[5] (.Q(
      mem_backbone_0_pmem_dout_bckup[5]), .QN(), .CK(mem_backbone_0_n_13), .D(
      pmem_dout[5]), .RN(mem_backbone_0_n_2));
  AOI22_X1_LVT mem_backbone_0_i_39_11 (.ZN(mem_backbone_0_n_39_6), .A1(
      mem_backbone_0_n_39_0), .A2(pmem_dout[5]), .B1(
      mem_backbone_0_pmem_dout_bckup_sel), .B2(mem_backbone_0_pmem_dout_bckup[5]));
  INV_X1_LVT mem_backbone_0_i_39_12 (.ZN(fe_mdb_in[5]), .A(mem_backbone_0_n_39_6));
  DFFR_X1_LVT \mem_backbone_0_pmem_dout_bckup_reg[4] (.Q(
      mem_backbone_0_pmem_dout_bckup[4]), .QN(), .CK(mem_backbone_0_n_13), .D(
      pmem_dout[4]), .RN(mem_backbone_0_n_2));
  AOI22_X1_LVT mem_backbone_0_i_39_9 (.ZN(mem_backbone_0_n_39_5), .A1(
      mem_backbone_0_n_39_0), .A2(pmem_dout[4]), .B1(
      mem_backbone_0_pmem_dout_bckup_sel), .B2(mem_backbone_0_pmem_dout_bckup[4]));
  INV_X1_LVT mem_backbone_0_i_39_10 (.ZN(fe_mdb_in[4]), .A(mem_backbone_0_n_39_5));
  DFFR_X1_LVT \mem_backbone_0_pmem_dout_bckup_reg[3] (.Q(
      mem_backbone_0_pmem_dout_bckup[3]), .QN(), .CK(mem_backbone_0_n_13), .D(
      pmem_dout[3]), .RN(mem_backbone_0_n_2));
  AOI22_X1_LVT mem_backbone_0_i_39_7 (.ZN(mem_backbone_0_n_39_4), .A1(
      mem_backbone_0_n_39_0), .A2(pmem_dout[3]), .B1(
      mem_backbone_0_pmem_dout_bckup_sel), .B2(mem_backbone_0_pmem_dout_bckup[3]));
  INV_X1_LVT mem_backbone_0_i_39_8 (.ZN(fe_mdb_in[3]), .A(mem_backbone_0_n_39_4));
  DFFR_X1_LVT \mem_backbone_0_pmem_dout_bckup_reg[2] (.Q(
      mem_backbone_0_pmem_dout_bckup[2]), .QN(), .CK(mem_backbone_0_n_13), .D(
      pmem_dout[2]), .RN(mem_backbone_0_n_2));
  AOI22_X1_LVT mem_backbone_0_i_39_5 (.ZN(mem_backbone_0_n_39_3), .A1(
      mem_backbone_0_n_39_0), .A2(pmem_dout[2]), .B1(
      mem_backbone_0_pmem_dout_bckup_sel), .B2(mem_backbone_0_pmem_dout_bckup[2]));
  INV_X1_LVT mem_backbone_0_i_39_6 (.ZN(fe_mdb_in[2]), .A(mem_backbone_0_n_39_3));
  DFFR_X1_LVT \mem_backbone_0_pmem_dout_bckup_reg[1] (.Q(
      mem_backbone_0_pmem_dout_bckup[1]), .QN(), .CK(mem_backbone_0_n_13), .D(
      pmem_dout[1]), .RN(mem_backbone_0_n_2));
  AOI22_X1_LVT mem_backbone_0_i_39_3 (.ZN(mem_backbone_0_n_39_2), .A1(
      mem_backbone_0_n_39_0), .A2(pmem_dout[1]), .B1(
      mem_backbone_0_pmem_dout_bckup_sel), .B2(mem_backbone_0_pmem_dout_bckup[1]));
  INV_X1_LVT mem_backbone_0_i_39_4 (.ZN(fe_mdb_in[1]), .A(mem_backbone_0_n_39_2));
  DFFR_X1_LVT \mem_backbone_0_pmem_dout_bckup_reg[0] (.Q(
      mem_backbone_0_pmem_dout_bckup[0]), .QN(), .CK(mem_backbone_0_n_13), .D(
      pmem_dout[0]), .RN(mem_backbone_0_n_2));
  AOI22_X1_LVT mem_backbone_0_i_39_1 (.ZN(mem_backbone_0_n_39_1), .A1(
      mem_backbone_0_n_39_0), .A2(pmem_dout[0]), .B1(
      mem_backbone_0_pmem_dout_bckup[0]), .B2(mem_backbone_0_pmem_dout_bckup_sel));
  INV_X1_LVT mem_backbone_0_i_39_2 (.ZN(fe_mdb_in[0]), .A(mem_backbone_0_n_39_1));
  AND2_X1_LVT mem_backbone_0_i_40_0 (.ZN(fe_pmem_wait), .A1(
      mem_backbone_0_fe_pmem_en), .A2(mem_backbone_0_eu_pmem_en));
  INV_X1_LVT mem_backbone_0_i_41_0 (.ZN(mem_backbone_0_n_16), .A(dbg_mem_en));
  NAND2_X1_LVT mem_backbone_0_i_42_0 (.ZN(mem_backbone_0_n_42_0), .A1(
      mem_backbone_0_n_16), .A2(dma_en));
  NOR4_X1_LVT mem_backbone_0_i_42_1 (.ZN(dma_resp), .A1(mem_backbone_0_n_42_0), 
      .A2(mem_backbone_0_ext_dmem_sel), .A3(mem_backbone_0_ext_per_sel), .A4(
      mem_backbone_0_ext_pmem_sel));
  OR4_X1_LVT mem_backbone_0_i_43_0 (.ZN(mem_backbone_0_n_43_0), .A1(
      mem_backbone_0_ext_dmem_en), .A2(dma_resp), .A3(mem_backbone_0_ext_per_en), 
      .A4(mem_backbone_0_ext_pmem_en));
  AND2_X1_LVT mem_backbone_0_i_43_1 (.ZN(dma_ready), .A1(mem_backbone_0_n_43_0), 
      .A2(mem_backbone_0_n_16));
  DFFR_X1_LVT mem_backbone_0_dma_ready_dly_reg (.Q(mem_backbone_0_dma_ready_dly), 
      .QN(), .CK(mclk), .D(dma_ready), .RN(mem_backbone_0_n_2));
  AND2_X1_LVT mem_backbone_0_i_44_15 (.ZN(dma_dout[15]), .A1(
      mem_backbone_0_dma_ready_dly), .A2(dbg_mem_din[15]));
  AND2_X1_LVT mem_backbone_0_i_44_14 (.ZN(dma_dout[14]), .A1(
      mem_backbone_0_dma_ready_dly), .A2(dbg_mem_din[14]));
  AND2_X1_LVT mem_backbone_0_i_44_13 (.ZN(dma_dout[13]), .A1(
      mem_backbone_0_dma_ready_dly), .A2(dbg_mem_din[13]));
  AND2_X1_LVT mem_backbone_0_i_44_12 (.ZN(dma_dout[12]), .A1(
      mem_backbone_0_dma_ready_dly), .A2(dbg_mem_din[12]));
  AND2_X1_LVT mem_backbone_0_i_44_11 (.ZN(dma_dout[11]), .A1(
      mem_backbone_0_dma_ready_dly), .A2(dbg_mem_din[11]));
  AND2_X1_LVT mem_backbone_0_i_44_10 (.ZN(dma_dout[10]), .A1(
      mem_backbone_0_dma_ready_dly), .A2(dbg_mem_din[10]));
  AND2_X1_LVT mem_backbone_0_i_44_9 (.ZN(dma_dout[9]), .A1(
      mem_backbone_0_dma_ready_dly), .A2(dbg_mem_din[9]));
  AND2_X1_LVT mem_backbone_0_i_44_8 (.ZN(dma_dout[8]), .A1(
      mem_backbone_0_dma_ready_dly), .A2(dbg_mem_din[8]));
  AND2_X1_LVT mem_backbone_0_i_44_7 (.ZN(dma_dout[7]), .A1(
      mem_backbone_0_dma_ready_dly), .A2(dbg_mem_din[7]));
  AND2_X1_LVT mem_backbone_0_i_44_6 (.ZN(dma_dout[6]), .A1(
      mem_backbone_0_dma_ready_dly), .A2(dbg_mem_din[6]));
  AND2_X1_LVT mem_backbone_0_i_44_5 (.ZN(dma_dout[5]), .A1(
      mem_backbone_0_dma_ready_dly), .A2(dbg_mem_din[5]));
  AND2_X1_LVT mem_backbone_0_i_44_4 (.ZN(dma_dout[4]), .A1(
      mem_backbone_0_dma_ready_dly), .A2(dbg_mem_din[4]));
  AND2_X1_LVT mem_backbone_0_i_44_3 (.ZN(dma_dout[3]), .A1(
      mem_backbone_0_dma_ready_dly), .A2(dbg_mem_din[3]));
  AND2_X1_LVT mem_backbone_0_i_44_2 (.ZN(dma_dout[2]), .A1(
      mem_backbone_0_dma_ready_dly), .A2(dbg_mem_din[2]));
  AND2_X1_LVT mem_backbone_0_i_44_1 (.ZN(dma_dout[1]), .A1(
      mem_backbone_0_dma_ready_dly), .A2(dbg_mem_din[1]));
  AND2_X1_LVT mem_backbone_0_i_44_0 (.ZN(dma_dout[0]), .A1(dbg_mem_din[0]), .A2(
      mem_backbone_0_dma_ready_dly));
  INV_X1_LVT mem_backbone_0_i_45_0 (.ZN(mem_backbone_0_n_45_0), .A(
      mem_backbone_0_ext_per_en));
  AOI22_X1_LVT mem_backbone_0_i_45_15 (.ZN(mem_backbone_0_n_45_8), .A1(
      mem_backbone_0_n_45_0), .A2(eu_mab[8]), .B1(mem_backbone_0_ext_per_en), 
      .B2(mem_backbone_0_ext_mem_addr[7]));
  INV_X1_LVT mem_backbone_0_i_45_16 (.ZN(per_addr[7]), .A(mem_backbone_0_n_45_8));
  AOI22_X1_LVT mem_backbone_0_i_45_13 (.ZN(mem_backbone_0_n_45_7), .A1(
      mem_backbone_0_n_45_0), .A2(eu_mab[7]), .B1(mem_backbone_0_ext_per_en), 
      .B2(mem_backbone_0_ext_mem_addr[6]));
  INV_X1_LVT mem_backbone_0_i_45_14 (.ZN(per_addr[6]), .A(mem_backbone_0_n_45_7));
  AOI22_X1_LVT mem_backbone_0_i_45_11 (.ZN(mem_backbone_0_n_45_6), .A1(
      mem_backbone_0_n_45_0), .A2(eu_mab[6]), .B1(mem_backbone_0_ext_per_en), 
      .B2(mem_backbone_0_ext_mem_addr[5]));
  INV_X1_LVT mem_backbone_0_i_45_12 (.ZN(per_addr[5]), .A(mem_backbone_0_n_45_6));
  AOI22_X1_LVT mem_backbone_0_i_45_9 (.ZN(mem_backbone_0_n_45_5), .A1(
      mem_backbone_0_n_45_0), .A2(eu_mab[5]), .B1(mem_backbone_0_ext_per_en), 
      .B2(mem_backbone_0_ext_mem_addr[4]));
  INV_X1_LVT mem_backbone_0_i_45_10 (.ZN(per_addr[4]), .A(mem_backbone_0_n_45_5));
  AOI22_X1_LVT mem_backbone_0_i_45_7 (.ZN(mem_backbone_0_n_45_4), .A1(
      mem_backbone_0_n_45_0), .A2(eu_mab[4]), .B1(mem_backbone_0_ext_per_en), 
      .B2(mem_backbone_0_ext_mem_addr[3]));
  INV_X1_LVT mem_backbone_0_i_45_8 (.ZN(per_addr[3]), .A(mem_backbone_0_n_45_4));
  AOI22_X1_LVT mem_backbone_0_i_45_5 (.ZN(mem_backbone_0_n_45_3), .A1(
      mem_backbone_0_n_45_0), .A2(eu_mab[3]), .B1(mem_backbone_0_ext_per_en), 
      .B2(mem_backbone_0_ext_mem_addr[2]));
  INV_X1_LVT mem_backbone_0_i_45_6 (.ZN(per_addr[2]), .A(mem_backbone_0_n_45_3));
  AOI22_X1_LVT mem_backbone_0_i_45_3 (.ZN(mem_backbone_0_n_45_2), .A1(
      mem_backbone_0_n_45_0), .A2(eu_mab[2]), .B1(mem_backbone_0_ext_per_en), 
      .B2(mem_backbone_0_ext_mem_addr[1]));
  INV_X1_LVT mem_backbone_0_i_45_4 (.ZN(per_addr[1]), .A(mem_backbone_0_n_45_2));
  AOI22_X1_LVT mem_backbone_0_i_45_1 (.ZN(mem_backbone_0_n_45_1), .A1(
      mem_backbone_0_n_45_0), .A2(eu_mab[1]), .B1(mem_backbone_0_ext_mem_addr[0]), 
      .B2(mem_backbone_0_ext_per_en));
  INV_X1_LVT mem_backbone_0_i_45_2 (.ZN(per_addr[0]), .A(mem_backbone_0_n_45_1));
  INV_X1_LVT mem_backbone_0_i_46_0 (.ZN(mem_backbone_0_n_46_0), .A(
      mem_backbone_0_ext_per_en));
  AOI22_X1_LVT mem_backbone_0_i_46_31 (.ZN(mem_backbone_0_n_46_16), .A1(
      mem_backbone_0_n_46_0), .A2(eu_mdb_out[15]), .B1(mem_backbone_0_ext_per_en), 
      .B2(pmem_din[15]));
  INV_X1_LVT mem_backbone_0_i_46_32 (.ZN(per_din[15]), .A(mem_backbone_0_n_46_16));
  AOI22_X1_LVT mem_backbone_0_i_46_29 (.ZN(mem_backbone_0_n_46_15), .A1(
      mem_backbone_0_n_46_0), .A2(eu_mdb_out[14]), .B1(mem_backbone_0_ext_per_en), 
      .B2(pmem_din[14]));
  INV_X1_LVT mem_backbone_0_i_46_30 (.ZN(per_din[14]), .A(mem_backbone_0_n_46_15));
  AOI22_X1_LVT mem_backbone_0_i_46_27 (.ZN(mem_backbone_0_n_46_14), .A1(
      mem_backbone_0_n_46_0), .A2(eu_mdb_out[13]), .B1(mem_backbone_0_ext_per_en), 
      .B2(pmem_din[13]));
  INV_X1_LVT mem_backbone_0_i_46_28 (.ZN(per_din[13]), .A(mem_backbone_0_n_46_14));
  AOI22_X1_LVT mem_backbone_0_i_46_25 (.ZN(mem_backbone_0_n_46_13), .A1(
      mem_backbone_0_n_46_0), .A2(eu_mdb_out[12]), .B1(mem_backbone_0_ext_per_en), 
      .B2(pmem_din[12]));
  INV_X1_LVT mem_backbone_0_i_46_26 (.ZN(per_din[12]), .A(mem_backbone_0_n_46_13));
  AOI22_X1_LVT mem_backbone_0_i_46_23 (.ZN(mem_backbone_0_n_46_12), .A1(
      mem_backbone_0_n_46_0), .A2(eu_mdb_out[11]), .B1(mem_backbone_0_ext_per_en), 
      .B2(pmem_din[11]));
  INV_X1_LVT mem_backbone_0_i_46_24 (.ZN(per_din[11]), .A(mem_backbone_0_n_46_12));
  AOI22_X1_LVT mem_backbone_0_i_46_21 (.ZN(mem_backbone_0_n_46_11), .A1(
      mem_backbone_0_n_46_0), .A2(eu_mdb_out[10]), .B1(mem_backbone_0_ext_per_en), 
      .B2(pmem_din[10]));
  INV_X1_LVT mem_backbone_0_i_46_22 (.ZN(per_din[10]), .A(mem_backbone_0_n_46_11));
  AOI22_X1_LVT mem_backbone_0_i_46_19 (.ZN(mem_backbone_0_n_46_10), .A1(
      mem_backbone_0_n_46_0), .A2(eu_mdb_out[9]), .B1(mem_backbone_0_ext_per_en), 
      .B2(pmem_din[9]));
  INV_X1_LVT mem_backbone_0_i_46_20 (.ZN(per_din[9]), .A(mem_backbone_0_n_46_10));
  AOI22_X1_LVT mem_backbone_0_i_46_17 (.ZN(mem_backbone_0_n_46_9), .A1(
      mem_backbone_0_n_46_0), .A2(eu_mdb_out[8]), .B1(mem_backbone_0_ext_per_en), 
      .B2(pmem_din[8]));
  INV_X1_LVT mem_backbone_0_i_46_18 (.ZN(per_din[8]), .A(mem_backbone_0_n_46_9));
  AOI22_X1_LVT mem_backbone_0_i_46_15 (.ZN(mem_backbone_0_n_46_8), .A1(
      mem_backbone_0_n_46_0), .A2(eu_mdb_out[7]), .B1(mem_backbone_0_ext_per_en), 
      .B2(pmem_din[7]));
  INV_X1_LVT mem_backbone_0_i_46_16 (.ZN(per_din[7]), .A(mem_backbone_0_n_46_8));
  AOI22_X1_LVT mem_backbone_0_i_46_13 (.ZN(mem_backbone_0_n_46_7), .A1(
      mem_backbone_0_n_46_0), .A2(eu_mdb_out[6]), .B1(mem_backbone_0_ext_per_en), 
      .B2(pmem_din[6]));
  INV_X1_LVT mem_backbone_0_i_46_14 (.ZN(per_din[6]), .A(mem_backbone_0_n_46_7));
  AOI22_X1_LVT mem_backbone_0_i_46_11 (.ZN(mem_backbone_0_n_46_6), .A1(
      mem_backbone_0_n_46_0), .A2(eu_mdb_out[5]), .B1(mem_backbone_0_ext_per_en), 
      .B2(pmem_din[5]));
  INV_X1_LVT mem_backbone_0_i_46_12 (.ZN(per_din[5]), .A(mem_backbone_0_n_46_6));
  AOI22_X1_LVT mem_backbone_0_i_46_9 (.ZN(mem_backbone_0_n_46_5), .A1(
      mem_backbone_0_n_46_0), .A2(eu_mdb_out[4]), .B1(mem_backbone_0_ext_per_en), 
      .B2(pmem_din[4]));
  INV_X1_LVT mem_backbone_0_i_46_10 (.ZN(per_din[4]), .A(mem_backbone_0_n_46_5));
  AOI22_X1_LVT mem_backbone_0_i_46_7 (.ZN(mem_backbone_0_n_46_4), .A1(
      mem_backbone_0_n_46_0), .A2(eu_mdb_out[3]), .B1(mem_backbone_0_ext_per_en), 
      .B2(pmem_din[3]));
  INV_X1_LVT mem_backbone_0_i_46_8 (.ZN(per_din[3]), .A(mem_backbone_0_n_46_4));
  AOI22_X1_LVT mem_backbone_0_i_46_5 (.ZN(mem_backbone_0_n_46_3), .A1(
      mem_backbone_0_n_46_0), .A2(eu_mdb_out[2]), .B1(mem_backbone_0_ext_per_en), 
      .B2(pmem_din[2]));
  INV_X1_LVT mem_backbone_0_i_46_6 (.ZN(per_din[2]), .A(mem_backbone_0_n_46_3));
  AOI22_X1_LVT mem_backbone_0_i_46_3 (.ZN(mem_backbone_0_n_46_2), .A1(
      mem_backbone_0_n_46_0), .A2(eu_mdb_out[1]), .B1(mem_backbone_0_ext_per_en), 
      .B2(pmem_din[1]));
  INV_X1_LVT mem_backbone_0_i_46_4 (.ZN(per_din[1]), .A(mem_backbone_0_n_46_2));
  AOI22_X1_LVT mem_backbone_0_i_46_1 (.ZN(mem_backbone_0_n_46_1), .A1(
      mem_backbone_0_n_46_0), .A2(eu_mdb_out[0]), .B1(pmem_din[0]), .B2(
      mem_backbone_0_ext_per_en));
  INV_X1_LVT mem_backbone_0_i_46_2 (.ZN(per_din[0]), .A(mem_backbone_0_n_46_1));
  INV_X1_LVT mem_backbone_0_i_47_0 (.ZN(mem_backbone_0_n_47_0), .A(
      mem_backbone_0_ext_per_en));
  AOI22_X1_LVT mem_backbone_0_i_47_3 (.ZN(mem_backbone_0_n_47_2), .A1(
      mem_backbone_0_n_47_0), .A2(eu_mb_wr[1]), .B1(mem_backbone_0_ext_per_en), 
      .B2(mem_backbone_0_ext_mem_wr[1]));
  INV_X1_LVT mem_backbone_0_i_47_4 (.ZN(per_we[1]), .A(mem_backbone_0_n_47_2));
  AOI22_X1_LVT mem_backbone_0_i_47_1 (.ZN(mem_backbone_0_n_47_1), .A1(
      mem_backbone_0_n_47_0), .A2(eu_mb_wr[0]), .B1(mem_backbone_0_ext_mem_wr[0]), 
      .B2(mem_backbone_0_ext_per_en));
  INV_X1_LVT mem_backbone_0_i_47_2 (.ZN(per_we[0]), .A(mem_backbone_0_n_47_1));
  OR2_X1_LVT mem_backbone_0_i_48_0 (.ZN(per_en), .A1(mem_backbone_0_ext_per_en), 
      .A2(mem_backbone_0_eu_per_en));
  NOR2_X1_LVT mem_backbone_0_i_49_0 (.ZN(mem_backbone_0_n_49_0), .A1(
      mem_backbone_0_eu_pmem_en), .A2(mem_backbone_0_ext_pmem_en));
  AOI222_X1_LVT mem_backbone_0_i_49_21 (.ZN(mem_backbone_0_n_49_11), .A1(
      mem_backbone_0_n_49_0), .A2(n_10), .B1(mem_backbone_0_ext_pmem_en), .B2(
      mem_backbone_0_ext_mem_addr[10]), .C1(mem_backbone_0_eu_pmem_en), .C2(
      eu_mab[11]));
  INV_X1_LVT mem_backbone_0_i_49_22 (.ZN(pmem_addr[10]), .A(
      mem_backbone_0_n_49_11));
  AOI222_X1_LVT mem_backbone_0_i_49_19 (.ZN(mem_backbone_0_n_49_10), .A1(
      mem_backbone_0_n_49_0), .A2(n_9), .B1(mem_backbone_0_ext_pmem_en), .B2(
      mem_backbone_0_ext_mem_addr[9]), .C1(mem_backbone_0_eu_pmem_en), .C2(
      eu_mab[10]));
  INV_X1_LVT mem_backbone_0_i_49_20 (.ZN(pmem_addr[9]), .A(
      mem_backbone_0_n_49_10));
  AOI222_X1_LVT mem_backbone_0_i_49_17 (.ZN(mem_backbone_0_n_49_9), .A1(
      mem_backbone_0_n_49_0), .A2(n_8), .B1(mem_backbone_0_ext_pmem_en), .B2(
      mem_backbone_0_ext_mem_addr[8]), .C1(mem_backbone_0_eu_pmem_en), .C2(
      eu_mab[9]));
  INV_X1_LVT mem_backbone_0_i_49_18 (.ZN(pmem_addr[8]), .A(mem_backbone_0_n_49_9));
  AOI222_X1_LVT mem_backbone_0_i_49_15 (.ZN(mem_backbone_0_n_49_8), .A1(
      mem_backbone_0_n_49_0), .A2(n_7), .B1(mem_backbone_0_ext_pmem_en), .B2(
      mem_backbone_0_ext_mem_addr[7]), .C1(mem_backbone_0_eu_pmem_en), .C2(
      eu_mab[8]));
  INV_X1_LVT mem_backbone_0_i_49_16 (.ZN(pmem_addr[7]), .A(mem_backbone_0_n_49_8));
  AOI222_X1_LVT mem_backbone_0_i_49_13 (.ZN(mem_backbone_0_n_49_7), .A1(
      mem_backbone_0_n_49_0), .A2(n_6), .B1(mem_backbone_0_ext_pmem_en), .B2(
      mem_backbone_0_ext_mem_addr[6]), .C1(mem_backbone_0_eu_pmem_en), .C2(
      eu_mab[7]));
  INV_X1_LVT mem_backbone_0_i_49_14 (.ZN(pmem_addr[6]), .A(mem_backbone_0_n_49_7));
  AOI222_X1_LVT mem_backbone_0_i_49_11 (.ZN(mem_backbone_0_n_49_6), .A1(
      mem_backbone_0_n_49_0), .A2(n_5), .B1(mem_backbone_0_ext_pmem_en), .B2(
      mem_backbone_0_ext_mem_addr[5]), .C1(mem_backbone_0_eu_pmem_en), .C2(
      eu_mab[6]));
  INV_X1_LVT mem_backbone_0_i_49_12 (.ZN(pmem_addr[5]), .A(mem_backbone_0_n_49_6));
  AOI222_X1_LVT mem_backbone_0_i_49_9 (.ZN(mem_backbone_0_n_49_5), .A1(
      mem_backbone_0_n_49_0), .A2(n_4), .B1(mem_backbone_0_ext_pmem_en), .B2(
      mem_backbone_0_ext_mem_addr[4]), .C1(mem_backbone_0_eu_pmem_en), .C2(
      eu_mab[5]));
  INV_X1_LVT mem_backbone_0_i_49_10 (.ZN(pmem_addr[4]), .A(mem_backbone_0_n_49_5));
  AOI222_X1_LVT mem_backbone_0_i_49_7 (.ZN(mem_backbone_0_n_49_4), .A1(
      mem_backbone_0_n_49_0), .A2(n_3), .B1(mem_backbone_0_ext_pmem_en), .B2(
      mem_backbone_0_ext_mem_addr[3]), .C1(mem_backbone_0_eu_pmem_en), .C2(
      eu_mab[4]));
  INV_X1_LVT mem_backbone_0_i_49_8 (.ZN(pmem_addr[3]), .A(mem_backbone_0_n_49_4));
  AOI222_X1_LVT mem_backbone_0_i_49_5 (.ZN(mem_backbone_0_n_49_3), .A1(
      mem_backbone_0_n_49_0), .A2(n_2), .B1(mem_backbone_0_ext_pmem_en), .B2(
      mem_backbone_0_ext_mem_addr[2]), .C1(mem_backbone_0_eu_pmem_en), .C2(
      eu_mab[3]));
  INV_X1_LVT mem_backbone_0_i_49_6 (.ZN(pmem_addr[2]), .A(mem_backbone_0_n_49_3));
  AOI222_X1_LVT mem_backbone_0_i_49_3 (.ZN(mem_backbone_0_n_49_2), .A1(
      mem_backbone_0_n_49_0), .A2(n_1), .B1(mem_backbone_0_ext_pmem_en), .B2(
      mem_backbone_0_ext_mem_addr[1]), .C1(mem_backbone_0_eu_pmem_en), .C2(
      eu_mab[2]));
  INV_X1_LVT mem_backbone_0_i_49_4 (.ZN(pmem_addr[1]), .A(mem_backbone_0_n_49_2));
  AOI222_X1_LVT mem_backbone_0_i_49_1 (.ZN(mem_backbone_0_n_49_1), .A1(
      mem_backbone_0_n_49_0), .A2(n_0), .B1(mem_backbone_0_ext_mem_addr[0]), .B2(
      mem_backbone_0_ext_pmem_en), .C1(eu_mab[1]), .C2(mem_backbone_0_eu_pmem_en));
  INV_X1_LVT mem_backbone_0_i_49_2 (.ZN(pmem_addr[0]), .A(mem_backbone_0_n_49_1));
  NOR3_X1_LVT mem_backbone_0_i_50_0 (.ZN(pmem_cen), .A1(
      mem_backbone_0_fe_pmem_en), .A2(mem_backbone_0_ext_pmem_en), .A3(
      mem_backbone_0_eu_pmem_en));
  NAND2_X1_LVT mem_backbone_0_i_51_2 (.ZN(mem_backbone_0_n_51_1), .A1(
      mem_backbone_0_ext_pmem_en), .A2(mem_backbone_0_n_10));
  NAND2_X1_LVT mem_backbone_0_i_51_3 (.ZN(pmem_wen[1]), .A1(
      mem_backbone_0_n_51_1), .A2(mem_backbone_0_ext_pmem_en));
  NAND2_X1_LVT mem_backbone_0_i_51_0 (.ZN(mem_backbone_0_n_51_0), .A1(
      mem_backbone_0_n_9), .A2(mem_backbone_0_ext_pmem_en));
  NAND2_X1_LVT mem_backbone_0_i_51_1 (.ZN(pmem_wen[0]), .A1(mem_backbone_0_n_51_0), 
      .A2(mem_backbone_0_ext_pmem_en));
  INV_X1_LVT frontend_0_i_78_0 (.ZN(frontend_0_n_91), .A(puc_rst));
  DFFR_X1_LVT \frontend_0_i_state_reg[0] (.Q(frontend_0_i_state[0]), .QN(), .CK(
      cpu_mclk), .D(frontend_0_i_state_nxt_reg[0]), .RN(frontend_0_n_91));
  INV_X1_LVT frontend_0_i_76_2 (.ZN(frontend_0_n_76_2), .A(frontend_0_i_state[0]));
  INV_X1_LVT frontend_0_i_76_1 (.ZN(frontend_0_n_76_1), .A(frontend_0_i_state[2]));
  NOR3_X1_LVT frontend_0_i_76_3 (.ZN(frontend_0_n_76_3), .A1(frontend_0_n_76_1), 
      .A2(frontend_0_n_76_2), .A3(frontend_0_i_state[1]));
  INV_X1_LVT frontend_0_i_0_0 (.ZN(frontend_0_n_0_0), .A(cpu_halt_cmd));
  NAND2_X1_LVT frontend_0_i_0_1 (.ZN(frontend_0_cpu_halt_req), .A1(
      frontend_0_n_0_0), .A2(cpu_en_s));
  INV_X1_LVT frontend_0_i_1_0 (.ZN(frontend_0_n_0), .A(frontend_0_cpu_halt_req));
  INV_X1_LVT frontend_0_i_74_0 (.ZN(frontend_0_n_74_0), .A(frontend_0_n_0));
  NOR2_X1_LVT frontend_0_i_74_1 (.ZN(frontend_0_n_87), .A1(frontend_0_n_74_0), 
      .A2(cpuoff));
  INV_X1_LVT frontend_0_i_2_0 (.ZN(frontend_0_n_1), .A(cpu_halt_st));
  NAND2_X1_LVT frontend_0_i_4_0 (.ZN(frontend_0_n_4_0), .A1(frontend_0_n_1), .A2(
      frontend_0_n_0));
  NOR4_X1_LVT frontend_0_i_3_0 (.ZN(frontend_0_n_3_0), .A1(irq[10]), .A2(irq[11]), 
      .A3(irq[12]), .A4(irq[13]));
  NOR4_X1_LVT frontend_0_i_3_1 (.ZN(frontend_0_n_3_1), .A1(irq[2]), .A2(irq[3]), 
      .A3(irq[4]), .A4(irq[5]));
  NOR4_X1_LVT frontend_0_i_3_2 (.ZN(frontend_0_n_3_2), .A1(irq[6]), .A2(irq[7]), 
      .A3(irq[8]), .A4(irq[9]));
  NOR2_X1_LVT frontend_0_i_3_3 (.ZN(frontend_0_n_3_3), .A1(irq[0]), .A2(irq[1]));
  NAND4_X1_LVT frontend_0_i_3_4 (.ZN(frontend_0_n_2), .A1(frontend_0_n_3_0), .A2(
      frontend_0_n_3_1), .A3(frontend_0_n_3_2), .A4(frontend_0_n_3_3));
  OAI21_X1_LVT frontend_0_i_4_1 (.ZN(frontend_0_n_4_1), .A(gie), .B1(
      frontend_0_n_2), .B2(wdt_irq));
  INV_X1_LVT frontend_0_i_4_2 (.ZN(frontend_0_n_4_2), .A(nmi_pnd));
  AOI21_X1_LVT frontend_0_i_4_3 (.ZN(frontend_0_n_3), .A(frontend_0_n_4_0), .B1(
      frontend_0_n_4_1), .B2(frontend_0_n_4_2));
  AND2_X1_LVT frontend_0_i_74_2 (.ZN(frontend_0_n_88), .A1(frontend_0_n_0), .A2(
      frontend_0_n_3));
  NOR2_X1_LVT frontend_0_i_75_0 (.ZN(frontend_0_n_89), .A1(frontend_0_n_87), .A2(
      frontend_0_n_88));
  AND2_X1_LVT frontend_0_i_76_4 (.ZN(frontend_0_n_76_4), .A1(frontend_0_n_76_3), 
      .A2(frontend_0_n_89));
  INV_X1_LVT frontend_0_i_76_5 (.ZN(frontend_0_n_76_5), .A(frontend_0_i_state[1]));
  NOR3_X1_LVT frontend_0_i_76_6 (.ZN(frontend_0_n_76_6), .A1(frontend_0_n_76_5), 
      .A2(frontend_0_i_state[0]), .A3(frontend_0_i_state[2]));
  INV_X1_LVT frontend_0_i_55_0 (.ZN(frontend_0_n_55_0), .A(e_state[0]));
  INV_X1_LVT frontend_0_i_6_2 (.ZN(frontend_0_n_6_1), .A(frontend_0_i_state[2]));
  INV_X1_LVT frontend_0_i_6_3 (.ZN(frontend_0_n_6_2), .A(frontend_0_i_state[0]));
  NOR3_X1_LVT frontend_0_i_6_4 (.ZN(frontend_0_n_5), .A1(frontend_0_n_6_1), .A2(
      frontend_0_n_6_2), .A3(frontend_0_i_state[1]));
  OR2_X1_LVT frontend_0_i_49_2 (.ZN(frontend_0_n_55), .A1(frontend_0_n_5), .A2(
      frontend_0_cpu_halt_req));
  NOR3_X1_LVT frontend_0_i_8_0 (.ZN(frontend_0_n_10), .A1(fe_mdb_in[13]), .A2(
      fe_mdb_in[14]), .A3(fe_mdb_in[15]));
  NAND2_X1_LVT frontend_0_i_25_5 (.ZN(frontend_0_n_25_5), .A1(fe_mdb_in[7]), .A2(
      fe_mdb_in[8]));
  INV_X1_LVT frontend_0_i_25_6 (.ZN(frontend_0_n_25_6), .A(fe_mdb_in[9]));
  NOR2_X1_LVT frontend_0_i_25_14 (.ZN(frontend_0_n_29), .A1(frontend_0_n_25_5), 
      .A2(frontend_0_n_25_6));
  AND2_X1_LVT frontend_0_i_26_7 (.ZN(frontend_0_n_37), .A1(frontend_0_n_10), .A2(
      frontend_0_n_29));
  INV_X1_LVT frontend_0_i_27_8 (.ZN(frontend_0_n_27_1), .A(frontend_0_n_37));
  INV_X1_LVT frontend_0_i_25_0 (.ZN(frontend_0_n_25_0), .A(fe_mdb_in[7]));
  NAND2_X1_LVT frontend_0_i_25_4 (.ZN(frontend_0_n_25_4), .A1(frontend_0_n_25_0), 
      .A2(fe_mdb_in[8]));
  NOR2_X1_LVT frontend_0_i_25_13 (.ZN(frontend_0_n_28), .A1(frontend_0_n_25_4), 
      .A2(frontend_0_n_25_6));
  AND2_X1_LVT frontend_0_i_26_6 (.ZN(frontend_0_n_36), .A1(frontend_0_n_10), .A2(
      frontend_0_n_28));
  AND2_X1_LVT frontend_0_i_27_7 (.ZN(frontend_0_inst_so_nxt[6]), .A1(
      frontend_0_n_27_0), .A2(frontend_0_n_36));
  INV_X1_LVT frontend_0_i_7_0 (.ZN(frontend_0_n_9), .A(frontend_0_irq_detect));
  NAND2_X1_LVT frontend_0_i_11_0 (.ZN(frontend_0_n_11_0), .A1(fe_mdb_in[13]), 
      .A2(frontend_0_n_9));
  NOR3_X1_LVT frontend_0_i_11_1 (.ZN(frontend_0_inst_type_nxt), .A1(
      frontend_0_n_11_0), .A2(fe_mdb_in[14]), .A3(fe_mdb_in[15]));
  OR2_X1_LVT frontend_0_i_42_0 (.ZN(frontend_0_n_49), .A1(
      frontend_0_inst_so_nxt[6]), .A2(frontend_0_inst_type_nxt));
  INV_X1_LVT frontend_0_i_23_0 (.ZN(frontend_0_n_23_0), .A(fe_mdb_in[7]));
  NOR4_X1_LVT frontend_0_i_23_1 (.ZN(frontend_0_n_23_1), .A1(frontend_0_n_23_0), 
      .A2(fe_mdb_in[1]), .A3(fe_mdb_in[2]), .A4(fe_mdb_in[3]));
  INV_X1_LVT frontend_0_i_23_2 (.ZN(frontend_0_n_23_2), .A(fe_mdb_in[0]));
  NAND2_X1_LVT frontend_0_i_23_3 (.ZN(frontend_0_n_23_3), .A1(frontend_0_n_23_1), 
      .A2(frontend_0_n_23_2));
  NOR4_X1_LVT frontend_0_i_23_4 (.ZN(frontend_0_n_23_4), .A1(fe_mdb_in[0]), .A2(
      fe_mdb_in[1]), .A3(fe_mdb_in[2]), .A4(fe_mdb_in[3]));
  INV_X1_LVT frontend_0_i_23_5 (.ZN(frontend_0_n_23_5), .A(frontend_0_n_23_4));
  NAND2_X1_LVT frontend_0_i_23_6 (.ZN(frontend_0_n_23_6), .A1(frontend_0_n_23_3), 
      .A2(frontend_0_n_23_5));
  INV_X1_LVT frontend_0_i_23_7 (.ZN(frontend_0_n_23_7), .A(frontend_0_n_23_6));
  AOI22_X1_LVT frontend_0_i_23_8 (.ZN(frontend_0_n_23_8), .A1(frontend_0_n_23_3), 
      .A2(frontend_0_n_23_4), .B1(frontend_0_n_23_7), .B2(frontend_0_n_23_0));
  INV_X1_LVT frontend_0_i_23_9 (.ZN(frontend_0_n_23_9), .A(fe_mdb_in[2]));
  INV_X1_LVT frontend_0_i_23_10 (.ZN(frontend_0_n_23_10), .A(fe_mdb_in[3]));
  NAND4_X1_LVT frontend_0_i_23_11 (.ZN(frontend_0_n_23_11), .A1(
      frontend_0_n_23_9), .A2(frontend_0_n_23_10), .A3(fe_mdb_in[7]), .A4(
      fe_mdb_in[1]));
  OR2_X1_LVT frontend_0_i_23_12 (.ZN(frontend_0_n_23_12), .A1(frontend_0_n_23_11), 
      .A2(fe_mdb_in[0]));
  OAI21_X1_LVT frontend_0_i_22_0 (.ZN(frontend_0_n_22_0), .A(frontend_0_n_9), 
      .B1(fe_mdb_in[14]), .B2(fe_mdb_in[15]));
  INV_X1_LVT frontend_0_i_22_1 (.ZN(frontend_0_n_17), .A(frontend_0_n_22_0));
  NAND2_X1_LVT frontend_0_i_23_13 (.ZN(frontend_0_n_23_13), .A1(
      frontend_0_n_23_12), .A2(frontend_0_n_17));
  INV_X1_LVT frontend_0_i_23_14 (.ZN(frontend_0_n_23_14), .A(frontend_0_n_23_13));
  NAND4_X1_LVT frontend_0_i_23_15 (.ZN(frontend_0_n_23_15), .A1(
      frontend_0_n_23_2), .A2(frontend_0_n_23_9), .A3(frontend_0_n_23_10), .A4(
      fe_mdb_in[1]));
  NAND2_X1_LVT frontend_0_i_23_16 (.ZN(frontend_0_n_23_16), .A1(
      frontend_0_n_23_14), .A2(frontend_0_n_23_15));
  OAI22_X1_LVT frontend_0_i_23_17 (.ZN(frontend_0_n_18), .A1(frontend_0_n_23_8), 
      .A2(frontend_0_n_23_16), .B1(frontend_0_n_23_15), .B2(frontend_0_n_23_13));
  NOR4_X1_LVT frontend_0_i_41_0 (.ZN(frontend_0_n_48), .A1(fe_mdb_in[0]), .A2(
      fe_mdb_in[1]), .A3(fe_mdb_in[2]), .A4(fe_mdb_in[3]));
  AOI21_X1_LVT frontend_0_i_44_0 (.ZN(frontend_0_n_44_0), .A(frontend_0_n_49), 
      .B1(frontend_0_n_18), .B2(frontend_0_n_48));
  INV_X1_LVT frontend_0_i_6_0 (.ZN(frontend_0_n_6_0), .A(frontend_0_i_state[1]));
  NOR3_X1_LVT frontend_0_i_6_1 (.ZN(frontend_0_n_4), .A1(frontend_0_n_6_0), .A2(
      frontend_0_i_state[0]), .A3(frontend_0_i_state[2]));
  OR2_X1_LVT frontend_0_i_61_0 (.ZN(frontend_0_n_73), .A1(frontend_0_n_67), .A2(
      exec_done));
  AND2_X1_LVT frontend_0_i_62_0 (.ZN(decode_noirq), .A1(frontend_0_n_4), .A2(
      frontend_0_n_73));
  OR2_X1_LVT frontend_0_i_63_0 (.ZN(frontend_0_decode), .A1(decode_noirq), .A2(
      frontend_0_irq_detect));
  INV_X1_LVT frontend_0_i_44_1 (.ZN(frontend_0_n_44_1), .A(frontend_0_decode));
  NOR2_X1_LVT frontend_0_i_44_2 (.ZN(frontend_0_n_51), .A1(frontend_0_n_44_0), 
      .A2(frontend_0_n_44_1));
  INV_X1_LVT frontend_0_i_45_0 (.ZN(frontend_0_n_45_0), .A(frontend_0_n_51));
  NAND3_X1_LVT frontend_0_i_45_1 (.ZN(frontend_0_n_45_1), .A1(frontend_0_n_45_0), 
      .A2(e_state[2]), .A3(e_state[3]));
  NOR3_X1_LVT frontend_0_i_45_2 (.ZN(frontend_0_n_45_2), .A1(frontend_0_n_45_1), 
      .A2(e_state[0]), .A3(e_state[1]));
  OR2_X1_LVT frontend_0_i_45_3 (.ZN(frontend_0_n_52), .A1(frontend_0_n_45_2), 
      .A2(frontend_0_n_51));
  CLKGATETST_X1_LVT frontend_0_clk_gate_exec_jmp_reg (.GCK(frontend_0_n_50), .CK(
      cpu_mclk), .E(frontend_0_n_52), .SE(1'b0));
  DFFR_X1_LVT frontend_0_exec_jmp_reg (.Q(frontend_0_exec_jmp), .QN(), .CK(
      frontend_0_n_50), .D(frontend_0_n_51), .RN(frontend_0_n_91));
  NOR2_X1_LVT frontend_0_i_59_0 (.ZN(frontend_0_n_59_0), .A1(
      frontend_0_exec_dst_wr), .A2(frontend_0_exec_jmp));
  AND2_X1_LVT frontend_0_i_9_0 (.ZN(frontend_0_n_11), .A1(frontend_0_n_10), .A2(
      frontend_0_n_9));
  CLKGATETST_X1_LVT frontend_0_clk_gate_inst_type_reg (.GCK(frontend_0_n_43), 
      .CK(cpu_mclk), .E(frontend_0_decode), .SE(1'b0));
  DFFR_X1_LVT \frontend_0_inst_type_reg[0] (.Q(inst_type[0]), .QN(), .CK(
      frontend_0_n_43), .D(frontend_0_n_11), .RN(frontend_0_n_91));
  INV_X1_LVT frontend_0_i_58_4 (.ZN(frontend_0_n_58_3), .A(e_state[1]));
  INV_X1_LVT frontend_0_i_58_2 (.ZN(frontend_0_n_58_2), .A(e_state[2]));
  NOR4_X1_LVT frontend_0_i_58_5 (.ZN(frontend_0_n_68), .A1(frontend_0_n_58_3), 
      .A2(frontend_0_n_58_2), .A3(e_state[0]), .A4(e_state[3]));
  AND2_X1_LVT frontend_0_i_37_0 (.ZN(frontend_0_n_45), .A1(inst_type[0]), .A2(
      frontend_0_n_68));
  INV_X1_LVT frontend_0_i_58_1 (.ZN(frontend_0_n_58_1), .A(e_state[0]));
  NOR4_X1_LVT frontend_0_i_58_6 (.ZN(frontend_0_n_69), .A1(frontend_0_n_58_2), 
      .A2(frontend_0_n_58_1), .A3(frontend_0_n_58_3), .A4(e_state[3]));
  NOR4_X1_LVT frontend_0_i_58_7 (.ZN(frontend_0_n_70), .A1(frontend_0_n_58_3), 
      .A2(frontend_0_n_58_0), .A3(e_state[0]), .A4(e_state[2]));
  OR2_X1_LVT frontend_0_i_38_0 (.ZN(frontend_0_n_46), .A1(frontend_0_n_69), .A2(
      frontend_0_n_70));
  INV_X1_LVT frontend_0_i_39_1 (.ZN(frontend_0_n_39_1), .A(frontend_0_n_46));
  INV_X1_LVT frontend_0_i_39_0 (.ZN(frontend_0_n_39_0), .A(frontend_0_n_45));
  NAND2_X1_LVT frontend_0_i_39_2 (.ZN(frontend_0_n_47), .A1(frontend_0_n_39_1), 
      .A2(frontend_0_n_39_0));
  CLKGATETST_X1_LVT frontend_0_clk_gate_exec_src_wr_reg (.GCK(frontend_0_n_44), 
      .CK(cpu_mclk), .E(frontend_0_n_47), .SE(1'b0));
  DFFR_X1_LVT frontend_0_exec_src_wr_reg (.Q(frontend_0_exec_src_wr), .QN(), .CK(
      frontend_0_n_44), .D(frontend_0_n_45), .RN(frontend_0_n_91));
  NAND3_X1_LVT frontend_0_i_59_1 (.ZN(frontend_0_n_59_1), .A1(frontend_0_n_59_0), 
      .A2(frontend_0_exec_src_wr), .A3(frontend_0_n_69));
  INV_X1_LVT frontend_0_i_59_2 (.ZN(frontend_0_n_59_2), .A(
      frontend_0_exec_src_wr));
  NOR4_X1_LVT frontend_0_i_58_9 (.ZN(frontend_0_n_72), .A1(frontend_0_n_58_0), 
      .A2(frontend_0_n_58_1), .A3(frontend_0_n_58_3), .A4(e_state[2]));
  NAND3_X1_LVT frontend_0_i_59_3 (.ZN(frontend_0_n_59_3), .A1(frontend_0_n_59_0), 
      .A2(frontend_0_n_59_2), .A3(frontend_0_n_72));
  INV_X1_LVT frontend_0_i_59_4 (.ZN(frontend_0_n_59_4), .A(frontend_0_exec_jmp));
  NAND3_X1_LVT frontend_0_i_59_5 (.ZN(frontend_0_n_59_5), .A1(frontend_0_n_59_4), 
      .A2(frontend_0_exec_dst_wr), .A3(frontend_0_n_70));
  NOR4_X1_LVT frontend_0_i_58_8 (.ZN(frontend_0_n_71), .A1(frontend_0_n_58_2), 
      .A2(frontend_0_n_58_0), .A3(e_state[0]), .A4(e_state[1]));
  NAND2_X1_LVT frontend_0_i_59_6 (.ZN(frontend_0_n_59_6), .A1(frontend_0_n_71), 
      .A2(frontend_0_exec_jmp));
  NAND4_X1_LVT frontend_0_i_59_7 (.ZN(exec_done), .A1(frontend_0_n_59_1), .A2(
      frontend_0_n_59_3), .A3(frontend_0_n_59_5), .A4(frontend_0_n_59_6));
  OAI21_X1_LVT frontend_0_i_60_0 (.ZN(frontend_0_n_60_0), .A(frontend_0_n_3), 
      .B1(frontend_0_n_5), .B2(exec_done));
  INV_X1_LVT frontend_0_i_60_1 (.ZN(frontend_0_irq_detect), .A(frontend_0_n_60_0));
  INV_X1_LVT frontend_0_i_27_0 (.ZN(frontend_0_n_27_0), .A(frontend_0_irq_detect));
  NAND2_X1_LVT frontend_0_i_27_9 (.ZN(frontend_0_inst_so_nxt[7]), .A1(
      frontend_0_n_27_1), .A2(frontend_0_n_27_0));
  AND2_X1_LVT frontend_0_i_49_3 (.ZN(frontend_0_n_56), .A1(frontend_0_n_1), .A2(
      frontend_0_inst_so_nxt[7]));
  NOR2_X1_LVT frontend_0_i_50_0 (.ZN(frontend_0_n_50_0), .A1(frontend_0_n_55), 
      .A2(frontend_0_n_56));
  INV_X1_LVT frontend_0_i_50_1 (.ZN(frontend_0_n_50_1), .A(frontend_0_n_50_0));
  NOR2_X1_LVT frontend_0_i_50_2 (.ZN(frontend_0_n_50_2), .A1(frontend_0_n_50_1), 
      .A2(cpuoff));
  INV_X1_LVT frontend_0_i_50_3 (.ZN(frontend_0_n_50_3), .A(frontend_0_n_50_2));
  INV_X1_LVT frontend_0_i_10_0 (.ZN(frontend_0_n_10_0), .A(frontend_0_n_11));
  AOI22_X1_LVT frontend_0_i_10_1 (.ZN(frontend_0_n_10_1), .A1(frontend_0_n_10_0), 
      .A2(fe_mdb_in[8]), .B1(fe_mdb_in[0]), .B2(frontend_0_n_11));
  INV_X1_LVT frontend_0_i_10_2 (.ZN(frontend_0_src_reg[0]), .A(frontend_0_n_10_1));
  AOI22_X1_LVT frontend_0_i_10_3 (.ZN(frontend_0_n_10_2), .A1(frontend_0_n_10_0), 
      .A2(fe_mdb_in[9]), .B1(frontend_0_n_11), .B2(fe_mdb_in[1]));
  INV_X1_LVT frontend_0_i_10_4 (.ZN(frontend_0_src_reg[1]), .A(frontend_0_n_10_2));
  AOI22_X1_LVT frontend_0_i_10_5 (.ZN(frontend_0_n_10_3), .A1(frontend_0_n_10_0), 
      .A2(fe_mdb_in[10]), .B1(frontend_0_n_11), .B2(fe_mdb_in[2]));
  INV_X1_LVT frontend_0_i_10_6 (.ZN(frontend_0_src_reg[2]), .A(frontend_0_n_10_3));
  AOI22_X1_LVT frontend_0_i_10_7 (.ZN(frontend_0_n_10_4), .A1(frontend_0_n_10_0), 
      .A2(fe_mdb_in[11]), .B1(frontend_0_n_11), .B2(fe_mdb_in[3]));
  INV_X1_LVT frontend_0_i_10_8 (.ZN(frontend_0_src_reg[3]), .A(frontend_0_n_10_4));
  NOR4_X1_LVT frontend_0_i_12_12 (.ZN(frontend_0_n_12_11), .A1(
      frontend_0_src_reg[0]), .A2(frontend_0_src_reg[1]), .A3(
      frontend_0_src_reg[2]), .A4(frontend_0_src_reg[3]));
  INV_X1_LVT frontend_0_i_12_16 (.ZN(frontend_0_n_12_12), .A(frontend_0_n_12_11));
  INV_X1_LVT frontend_0_i_12_6 (.ZN(frontend_0_n_12_6), .A(frontend_0_src_reg[0]));
  INV_X1_LVT frontend_0_i_12_7 (.ZN(frontend_0_n_12_7), .A(frontend_0_src_reg[1]));
  NOR4_X1_LVT frontend_0_i_12_8 (.ZN(frontend_0_n_12_8), .A1(frontend_0_n_12_6), 
      .A2(frontend_0_n_12_7), .A3(frontend_0_src_reg[2]), .A4(
      frontend_0_src_reg[3]));
  OR2_X1_LVT frontend_0_i_12_9 (.ZN(frontend_0_n_12_9), .A1(frontend_0_n_12_8), 
      .A2(frontend_0_inst_type_nxt));
  NOR4_X1_LVT frontend_0_i_12_11 (.ZN(frontend_0_n_12_10), .A1(frontend_0_n_12_7), 
      .A2(frontend_0_src_reg[0]), .A3(frontend_0_src_reg[2]), .A4(
      frontend_0_src_reg[3]));
  INV_X1_LVT frontend_0_i_12_1 (.ZN(frontend_0_n_12_1), .A(fe_mdb_in[5]));
  NAND2_X1_LVT frontend_0_i_12_3 (.ZN(frontend_0_n_12_3), .A1(frontend_0_n_12_1), 
      .A2(fe_mdb_in[4]));
  NOR4_X1_LVT frontend_0_i_12_17 (.ZN(frontend_0_inst_as_nxt[4]), .A1(
      frontend_0_n_12_12), .A2(frontend_0_n_12_9), .A3(frontend_0_n_12_10), .A4(
      frontend_0_n_12_3));
  INV_X1_LVT frontend_0_i_12_19 (.ZN(frontend_0_n_12_13), .A(frontend_0_n_12_10));
  NOR3_X1_LVT frontend_0_i_12_20 (.ZN(frontend_0_inst_as_nxt[6]), .A1(
      frontend_0_n_12_13), .A2(frontend_0_n_12_9), .A3(frontend_0_n_12_3));
  NOR4_X1_LVT frontend_0_i_12_13 (.ZN(frontend_0_inst_as_nxt[1]), .A1(
      frontend_0_n_12_9), .A2(frontend_0_n_12_10), .A3(frontend_0_n_12_3), .A4(
      frontend_0_n_12_11));
  OR3_X1_LVT frontend_0_i_48_0 (.ZN(frontend_0_src_acalc_pre), .A1(
      frontend_0_inst_as_nxt[4]), .A2(frontend_0_inst_as_nxt[6]), .A3(
      frontend_0_inst_as_nxt[1]));
  NOR2_X1_LVT frontend_0_i_50_4 (.ZN(frontend_0_n_50_4), .A1(frontend_0_n_50_3), 
      .A2(frontend_0_src_acalc_pre));
  OR2_X1_LVT frontend_0_i_12_2 (.ZN(frontend_0_n_12_2), .A1(frontend_0_n_12_1), 
      .A2(fe_mdb_in[4]));
  NOR3_X1_LVT frontend_0_i_12_14 (.ZN(frontend_0_inst_as_nxt[2]), .A1(
      frontend_0_n_12_9), .A2(frontend_0_n_12_10), .A3(frontend_0_n_12_2));
  NAND2_X1_LVT frontend_0_i_12_4 (.ZN(frontend_0_n_12_4), .A1(fe_mdb_in[4]), .A2(
      fe_mdb_in[5]));
  NOR4_X1_LVT frontend_0_i_12_15 (.ZN(frontend_0_inst_as_nxt[3]), .A1(
      frontend_0_n_12_9), .A2(frontend_0_n_12_10), .A3(frontend_0_n_12_11), .A4(
      frontend_0_n_12_4));
  NOR4_X1_LVT frontend_0_i_12_18 (.ZN(frontend_0_inst_as_nxt[5]), .A1(
      frontend_0_n_12_12), .A2(frontend_0_n_12_9), .A3(frontend_0_n_12_10), .A4(
      frontend_0_n_12_4));
  OR4_X1_LVT frontend_0_i_49_1 (.ZN(frontend_0_n_54), .A1(
      frontend_0_inst_as_nxt[2]), .A2(frontend_0_inst_as_nxt[3]), .A3(
      frontend_0_inst_as_nxt[5]), .A4(frontend_0_inst_so_nxt[6]));
  INV_X1_LVT frontend_0_i_50_5 (.ZN(frontend_0_n_50_5), .A(frontend_0_n_54));
  NAND2_X1_LVT frontend_0_i_50_6 (.ZN(frontend_0_n_50_6), .A1(frontend_0_n_50_4), 
      .A2(frontend_0_n_50_5));
  NOR2_X1_LVT frontend_0_i_23_19 (.ZN(frontend_0_n_20), .A1(frontend_0_n_23_3), 
      .A2(frontend_0_n_23_16));
  NOR3_X1_LVT frontend_0_i_23_18 (.ZN(frontend_0_n_19), .A1(frontend_0_n_23_16), 
      .A2(frontend_0_n_23_6), .A3(frontend_0_n_23_0));
  INV_X1_LVT frontend_0_i_23_20 (.ZN(frontend_0_n_23_17), .A(frontend_0_n_17));
  NOR2_X1_LVT frontend_0_i_23_21 (.ZN(frontend_0_inst_ad_nxt), .A1(
      frontend_0_n_23_12), .A2(frontend_0_n_23_17));
  OR3_X1_LVT frontend_0_i_47_0 (.ZN(frontend_0_dst_acalc_pre), .A1(
      frontend_0_n_20), .A2(frontend_0_n_19), .A3(frontend_0_inst_ad_nxt));
  NOR2_X1_LVT frontend_0_i_50_7 (.ZN(frontend_0_n_50_7), .A1(frontend_0_n_50_6), 
      .A2(frontend_0_dst_acalc_pre));
  INV_X1_LVT frontend_0_i_25_1 (.ZN(frontend_0_n_25_1), .A(fe_mdb_in[8]));
  NAND2_X1_LVT frontend_0_i_25_2 (.ZN(frontend_0_n_25_2), .A1(frontend_0_n_25_0), 
      .A2(frontend_0_n_25_1));
  NOR2_X1_LVT frontend_0_i_25_11 (.ZN(frontend_0_n_26), .A1(frontend_0_n_25_2), 
      .A2(frontend_0_n_25_6));
  AND2_X1_LVT frontend_0_i_26_4 (.ZN(frontend_0_n_34), .A1(frontend_0_n_10), .A2(
      frontend_0_n_26));
  AND2_X1_LVT frontend_0_i_27_5 (.ZN(frontend_0_inst_so_nxt[4]), .A1(
      frontend_0_n_27_0), .A2(frontend_0_n_34));
  NAND2_X1_LVT frontend_0_i_25_3 (.ZN(frontend_0_n_25_3), .A1(fe_mdb_in[7]), .A2(
      frontend_0_n_25_1));
  NOR2_X1_LVT frontend_0_i_25_12 (.ZN(frontend_0_n_27), .A1(frontend_0_n_25_3), 
      .A2(frontend_0_n_25_6));
  AND2_X1_LVT frontend_0_i_26_5 (.ZN(frontend_0_n_35), .A1(frontend_0_n_10), .A2(
      frontend_0_n_27));
  AND2_X1_LVT frontend_0_i_27_6 (.ZN(frontend_0_inst_so_nxt[5]), .A1(
      frontend_0_n_27_0), .A2(frontend_0_n_35));
  OR2_X1_LVT frontend_0_i_49_0 (.ZN(frontend_0_n_53), .A1(
      frontend_0_inst_so_nxt[4]), .A2(frontend_0_inst_so_nxt[5]));
  INV_X1_LVT frontend_0_i_50_8 (.ZN(frontend_0_n_50_8), .A(frontend_0_n_53));
  NAND2_X1_LVT frontend_0_i_50_9 (.ZN(frontend_0_n_50_9), .A1(frontend_0_n_50_7), 
      .A2(frontend_0_n_50_8));
  NAND2_X1_LVT frontend_0_i_50_17 (.ZN(frontend_0_n_50_16), .A1(
      frontend_0_n_50_4), .A2(frontend_0_n_54));
  INV_X1_LVT frontend_0_i_50_12 (.ZN(frontend_0_n_50_12), .A(frontend_0_n_56));
  NAND3_X1_LVT frontend_0_i_50_18 (.ZN(frontend_0_n_58), .A1(frontend_0_n_50_9), 
      .A2(frontend_0_n_50_16), .A3(frontend_0_n_50_12));
  AND2_X1_LVT frontend_0_i_55_36 (.ZN(frontend_0_n_55_35), .A1(frontend_0_n_55_6), 
      .A2(frontend_0_n_58));
  NOR4_X1_LVT frontend_0_i_55_18 (.ZN(frontend_0_n_55_18), .A1(e_state[0]), .A2(
      e_state[1]), .A3(e_state[2]), .A4(e_state[3]));
  NAND4_X1_LVT frontend_0_i_55_23 (.ZN(frontend_0_n_55_23), .A1(
      frontend_0_n_55_1), .A2(frontend_0_n_55_10), .A3(e_state[0]), .A4(
      e_state[3]));
  INV_X1_LVT frontend_0_i_55_37 (.ZN(frontend_0_n_55_36), .A(frontend_0_n_55_23));
  NOR4_X1_LVT frontend_0_i_55_38 (.ZN(frontend_0_n_55_37), .A1(
      frontend_0_n_55_35), .A2(frontend_0_n_55_18), .A3(frontend_0_n_55_21), .A4(
      frontend_0_n_55_36));
  NOR4_X1_LVT frontend_0_i_55_30 (.ZN(frontend_0_n_55_30), .A1(frontend_0_n_55_0), 
      .A2(frontend_0_n_55_10), .A3(e_state[1]), .A4(e_state[3]));
  NOR3_X1_LVT frontend_0_i_6_5 (.ZN(frontend_0_n_6), .A1(frontend_0_n_6_0), .A2(
      frontend_0_n_6_2), .A3(frontend_0_i_state[2]));
  CLKGATETST_X1_LVT frontend_0_clk_gate_inst_as_reg (.GCK(frontend_0_n_12), .CK(
      cpu_mclk), .E(frontend_0_decode), .SE(1'b0));
  DFFR_X1_LVT \frontend_0_inst_as_reg[6] (.Q(inst_as[6]), .QN(), .CK(
      frontend_0_n_12), .D(frontend_0_inst_as_nxt[6]), .RN(frontend_0_n_91));
  DFFR_X1_LVT \frontend_0_inst_as_reg[1] (.Q(inst_as[1]), .QN(), .CK(
      frontend_0_n_12), .D(frontend_0_inst_as_nxt[1]), .RN(frontend_0_n_91));
  DFFR_X1_LVT \frontend_0_inst_as_reg[5] (.Q(inst_as[5]), .QN(), .CK(
      frontend_0_n_12), .D(frontend_0_inst_as_nxt[5]), .RN(frontend_0_n_91));
  DFFR_X1_LVT \frontend_0_inst_as_reg[4] (.Q(inst_as[4]), .QN(), .CK(
      frontend_0_n_12), .D(frontend_0_inst_as_nxt[4]), .RN(frontend_0_n_91));
  OR4_X1_LVT frontend_0_i_15_0 (.ZN(frontend_0_is_sext), .A1(inst_as[6]), .A2(
      inst_as[1]), .A3(inst_as[5]), .A4(inst_as[4]));
  AND2_X1_LVT frontend_0_i_30_0 (.ZN(frontend_0_inst_sext_rdy), .A1(
      frontend_0_n_6), .A2(frontend_0_is_sext));
  NAND2_X1_LVT frontend_0_i_55_39 (.ZN(frontend_0_n_55_38), .A1(
      frontend_0_n_55_30), .A2(frontend_0_inst_sext_rdy));
  INV_X1_LVT frontend_0_i_55_4 (.ZN(frontend_0_n_55_4), .A(e_state[3]));
  NAND4_X1_LVT frontend_0_i_55_32 (.ZN(frontend_0_n_55_32), .A1(
      frontend_0_n_55_0), .A2(frontend_0_n_55_4), .A3(e_state[1]), .A4(
      e_state[2]));
  INV_X1_LVT frontend_0_i_55_33 (.ZN(frontend_0_n_55_33), .A(frontend_0_n_55_32));
  CLKGATETST_X1_LVT frontend_0_clk_gate_inst_so_reg (.GCK(frontend_0_n_38), .CK(
      cpu_mclk), .E(frontend_0_decode), .SE(1'b0));
  DFFR_X1_LVT \frontend_0_inst_so_reg[6] (.Q(inst_so[6]), .QN(), .CK(
      frontend_0_n_38), .D(frontend_0_inst_so_nxt[6]), .RN(frontend_0_n_91));
  DFFR_X1_LVT \frontend_0_inst_so_reg[4] (.Q(inst_so[4]), .QN(), .CK(
      frontend_0_n_38), .D(frontend_0_inst_so_nxt[4]), .RN(frontend_0_n_91));
  DFFR_X1_LVT \frontend_0_inst_so_reg[5] (.Q(inst_so[5]), .QN(), .CK(
      frontend_0_n_38), .D(frontend_0_inst_so_nxt[5]), .RN(frontend_0_n_91));
  OR2_X1_LVT frontend_0_i_29_0 (.ZN(frontend_0_n_39), .A1(inst_so[4]), .A2(
      inst_so[5]));
  OR2_X1_LVT frontend_0_i_52_0 (.ZN(frontend_0_n_62), .A1(inst_so[6]), .A2(
      frontend_0_n_39));
  CLKGATETST_X1_LVT frontend_0_clk_gate_inst_ad_reg (.GCK(frontend_0_n_21), .CK(
      cpu_mclk), .E(frontend_0_decode), .SE(1'b0));
  DFFR_X1_LVT \frontend_0_inst_ad_reg[4] (.Q(inst_ad[4]), .QN(), .CK(
      frontend_0_n_21), .D(frontend_0_n_20), .RN(frontend_0_n_91));
  DFFR_X1_LVT \frontend_0_inst_ad_reg[1] (.Q(inst_ad[1]), .QN(), .CK(
      frontend_0_n_21), .D(frontend_0_n_19), .RN(frontend_0_n_91));
  DFFR_X1_LVT \frontend_0_inst_ad_reg[6] (.Q(inst_ad[6]), .QN(), .CK(
      frontend_0_n_21), .D(frontend_0_inst_ad_nxt), .RN(frontend_0_n_91));
  OR3_X1_LVT frontend_0_i_52_1 (.ZN(frontend_0_n_63), .A1(inst_ad[4]), .A2(
      inst_ad[1]), .A3(inst_ad[6]));
  NOR2_X1_LVT frontend_0_i_53_0 (.ZN(frontend_0_n_64), .A1(frontend_0_n_62), .A2(
      frontend_0_n_63));
  NAND2_X1_LVT frontend_0_i_55_40 (.ZN(frontend_0_n_55_39), .A1(
      frontend_0_n_55_33), .A2(frontend_0_n_64));
  NAND4_X1_LVT frontend_0_i_55_11 (.ZN(frontend_0_n_55_11), .A1(
      frontend_0_n_55_10), .A2(e_state[0]), .A3(e_state[1]), .A4(e_state[3]));
  INV_X1_LVT frontend_0_i_55_41 (.ZN(frontend_0_n_55_40), .A(frontend_0_n_55_11));
  NOR2_X1_LVT frontend_0_i_55_12 (.ZN(frontend_0_n_55_12), .A1(
      frontend_0_exec_jmp), .A2(frontend_0_exec_dst_wr));
  NAND2_X1_LVT frontend_0_i_55_16 (.ZN(frontend_0_n_55_16), .A1(
      frontend_0_n_55_12), .A2(frontend_0_exec_src_wr));
  INV_X1_LVT frontend_0_i_55_13 (.ZN(frontend_0_n_55_13), .A(frontend_0_n_55_12));
  NOR2_X1_LVT frontend_0_i_55_14 (.ZN(frontend_0_n_55_14), .A1(
      frontend_0_n_55_13), .A2(frontend_0_exec_src_wr));
  INV_X1_LVT frontend_0_i_55_43 (.ZN(frontend_0_n_55_42), .A(frontend_0_n_55_14));
  INV_X1_LVT frontend_0_i_55_44 (.ZN(frontend_0_n_55_43), .A(frontend_0_n_58));
  OAI211_X1_LVT frontend_0_i_55_45 (.ZN(frontend_0_n_55_44), .A(
      frontend_0_n_55_16), .B(frontend_0_n_55_41), .C1(frontend_0_n_55_42), .C2(
      frontend_0_n_55_43));
  NAND2_X1_LVT frontend_0_i_55_46 (.ZN(frontend_0_n_55_45), .A1(
      frontend_0_n_55_40), .A2(frontend_0_n_55_44));
  AND4_X1_LVT frontend_0_i_55_47 (.ZN(frontend_0_n_55_46), .A1(
      frontend_0_n_55_37), .A2(frontend_0_n_55_38), .A3(frontend_0_n_55_39), .A4(
      frontend_0_n_55_45));
  NAND4_X1_LVT frontend_0_i_55_26 (.ZN(frontend_0_n_55_26), .A1(
      frontend_0_n_55_0), .A2(frontend_0_n_55_10), .A3(e_state[1]), .A4(
      e_state[3]));
  INV_X1_LVT frontend_0_i_55_27 (.ZN(frontend_0_n_55_27), .A(frontend_0_n_55_26));
  INV_X1_LVT frontend_0_i_55_28 (.ZN(frontend_0_n_55_28), .A(frontend_0_exec_jmp));
  NAND3_X1_LVT frontend_0_i_55_48 (.ZN(frontend_0_n_55_47), .A1(
      frontend_0_n_55_27), .A2(frontend_0_n_55_28), .A3(frontend_0_n_58));
  NAND4_X1_LVT frontend_0_i_55_3 (.ZN(frontend_0_n_55_3), .A1(frontend_0_n_55_1), 
      .A2(e_state[0]), .A3(e_state[2]), .A4(e_state[3]));
  NAND4_X1_LVT frontend_0_i_55_5 (.ZN(frontend_0_n_55_5), .A1(frontend_0_n_55_4), 
      .A2(e_state[0]), .A3(e_state[1]), .A4(e_state[2]));
  AND4_X1_LVT frontend_0_i_55_49 (.ZN(frontend_0_n_55_48), .A1(
      frontend_0_n_55_26), .A2(frontend_0_n_55_3), .A3(frontend_0_n_55_11), .A4(
      frontend_0_n_55_5));
  NAND4_X1_LVT frontend_0_i_55_50 (.ZN(frontend_0_n_55_49), .A1(
      frontend_0_n_55_48), .A2(frontend_0_n_55_32), .A3(frontend_0_n_55_23), .A4(
      frontend_0_n_55_2));
  NOR4_X1_LVT frontend_0_i_55_8 (.ZN(frontend_0_n_55_8), .A1(frontend_0_n_55_4), 
      .A2(e_state[0]), .A3(e_state[1]), .A4(e_state[2]));
  NOR4_X1_LVT frontend_0_i_55_51 (.ZN(frontend_0_n_55_50), .A1(frontend_0_n_55_0), 
      .A2(frontend_0_n_55_1), .A3(e_state[2]), .A4(e_state[3]));
  NOR4_X1_LVT frontend_0_i_55_52 (.ZN(frontend_0_n_55_51), .A1(
      frontend_0_n_55_49), .A2(frontend_0_n_55_8), .A3(frontend_0_n_55_50), .A4(
      frontend_0_n_55_30));
  NAND4_X1_LVT frontend_0_i_55_20 (.ZN(frontend_0_n_55_20), .A1(
      frontend_0_n_55_0), .A2(frontend_0_n_55_10), .A3(frontend_0_n_55_4), .A4(
      e_state[1]));
  NAND4_X1_LVT frontend_0_i_55_53 (.ZN(frontend_0_n_55_52), .A1(
      frontend_0_n_55_1), .A2(frontend_0_n_55_10), .A3(frontend_0_n_55_4), .A4(
      e_state[0]));
  INV_X1_LVT frontend_0_i_55_22 (.ZN(frontend_0_n_55_22), .A(frontend_0_n_55_21));
  NAND4_X1_LVT frontend_0_i_55_54 (.ZN(frontend_0_n_55_53), .A1(
      frontend_0_n_55_51), .A2(frontend_0_n_55_20), .A3(frontend_0_n_55_52), .A4(
      frontend_0_n_55_22));
  OAI211_X1_LVT frontend_0_i_55_55 (.ZN(frontend_0_e_state_nxt_reg[1]), .A(
      frontend_0_n_55_46), .B(frontend_0_n_55_47), .C1(frontend_0_n_55_53), .C2(
      frontend_0_n_55_18));
  DFFR_X1_LVT \frontend_0_e_state_reg[1] (.Q(e_state[1]), .QN(), .CK(cpu_mclk), 
      .D(frontend_0_e_state_nxt_reg[1]), .RN(frontend_0_n_91));
  INV_X1_LVT frontend_0_i_55_1 (.ZN(frontend_0_n_55_1), .A(e_state[1]));
  NAND4_X1_LVT frontend_0_i_55_2 (.ZN(frontend_0_n_55_2), .A1(frontend_0_n_55_0), 
      .A2(frontend_0_n_55_1), .A3(e_state[2]), .A4(e_state[3]));
  NAND3_X1_LVT frontend_0_i_55_6 (.ZN(frontend_0_n_55_6), .A1(frontend_0_n_55_2), 
      .A2(frontend_0_n_55_3), .A3(frontend_0_n_55_5));
  NAND2_X1_LVT frontend_0_i_50_10 (.ZN(frontend_0_n_50_10), .A1(
      frontend_0_n_50_2), .A2(frontend_0_src_acalc_pre));
  NAND2_X1_LVT frontend_0_i_50_11 (.ZN(frontend_0_n_50_11), .A1(
      frontend_0_n_50_0), .A2(cpuoff));
  NAND2_X1_LVT frontend_0_i_50_13 (.ZN(frontend_0_n_50_13), .A1(
      frontend_0_n_50_12), .A2(frontend_0_n_55));
  AND4_X1_LVT frontend_0_i_50_14 (.ZN(frontend_0_n_50_14), .A1(frontend_0_n_50_9), 
      .A2(frontend_0_n_50_10), .A3(frontend_0_n_50_11), .A4(frontend_0_n_50_13));
  NAND2_X1_LVT frontend_0_i_50_15 (.ZN(frontend_0_n_50_15), .A1(
      frontend_0_n_50_7), .A2(frontend_0_n_53));
  NAND2_X1_LVT frontend_0_i_50_16 (.ZN(frontend_0_n_57), .A1(frontend_0_n_50_14), 
      .A2(frontend_0_n_50_15));
  AND2_X1_LVT frontend_0_i_55_7 (.ZN(frontend_0_n_55_7), .A1(frontend_0_n_55_6), 
      .A2(frontend_0_n_57));
  INV_X1_LVT frontend_0_i_16_0 (.ZN(frontend_0_n_16_0), .A(frontend_0_n_6));
  NOR2_X1_LVT frontend_0_i_16_1 (.ZN(frontend_0_n_13), .A1(frontend_0_n_16_0), 
      .A2(frontend_0_is_sext));
  NOR3_X1_LVT frontend_0_i_6_6 (.ZN(frontend_0_n_7), .A1(frontend_0_n_6_1), .A2(
      frontend_0_i_state[0]), .A3(frontend_0_i_state[1]));
  OR2_X1_LVT frontend_0_i_17_0 (.ZN(frontend_0_inst_dext_rdy), .A1(
      frontend_0_n_13), .A2(frontend_0_n_7));
  NAND2_X1_LVT frontend_0_i_19_0 (.ZN(frontend_0_n_19_0), .A1(e_state[0]), .A2(
      e_state[3]));
  OR3_X1_LVT frontend_0_i_19_1 (.ZN(frontend_0_n_19_1), .A1(frontend_0_n_19_0), 
      .A2(e_state[1]), .A3(e_state[2]));
  AND2_X1_LVT frontend_0_i_19_2 (.ZN(frontend_0_n_15), .A1(frontend_0_n_19_1), 
      .A2(frontend_0_inst_dext_rdy));
  INV_X1_LVT frontend_0_i_20_3 (.ZN(frontend_0_n_20_3), .A(
      frontend_0_inst_dext_rdy));
  NAND2_X1_LVT frontend_0_i_20_0 (.ZN(frontend_0_n_20_0), .A1(e_state[0]), .A2(
      e_state[3]));
  NOR3_X1_LVT frontend_0_i_20_1 (.ZN(frontend_0_n_20_1), .A1(frontend_0_n_20_0), 
      .A2(e_state[1]), .A3(e_state[2]));
  INV_X1_LVT frontend_0_i_20_2 (.ZN(frontend_0_n_20_2), .A(frontend_0_n_20_1));
  NAND2_X1_LVT frontend_0_i_20_4 (.ZN(frontend_0_n_16), .A1(frontend_0_n_20_3), 
      .A2(frontend_0_n_20_2));
  CLKGATETST_X1_LVT frontend_0_clk_gate_exec_dext_rdy_reg (.GCK(frontend_0_n_14), 
      .CK(cpu_mclk), .E(frontend_0_n_16), .SE(1'b0));
  DFFR_X1_LVT frontend_0_exec_dext_rdy_reg (.Q(frontend_0_exec_dext_rdy), .QN(), 
      .CK(frontend_0_n_14), .D(frontend_0_n_15), .RN(frontend_0_n_91));
  OR2_X1_LVT frontend_0_i_51_0 (.ZN(frontend_0_n_61), .A1(
      frontend_0_inst_dext_rdy), .A2(frontend_0_exec_dext_rdy));
  AND2_X1_LVT frontend_0_i_55_9 (.ZN(frontend_0_n_55_9), .A1(frontend_0_n_55_8), 
      .A2(frontend_0_n_61));
  NAND2_X1_LVT frontend_0_i_55_15 (.ZN(frontend_0_n_55_15), .A1(
      frontend_0_n_55_14), .A2(frontend_0_n_57));
  AOI21_X1_LVT frontend_0_i_55_17 (.ZN(frontend_0_n_55_17), .A(
      frontend_0_n_55_11), .B1(frontend_0_n_55_15), .B2(frontend_0_n_55_16));
  INV_X1_LVT frontend_0_i_55_19 (.ZN(frontend_0_n_55_19), .A(frontend_0_n_55_18));
  NAND4_X1_LVT frontend_0_i_55_24 (.ZN(frontend_0_n_55_24), .A1(
      frontend_0_n_55_19), .A2(frontend_0_n_55_20), .A3(frontend_0_n_55_22), .A4(
      frontend_0_n_55_23));
  NOR4_X1_LVT frontend_0_i_55_25 (.ZN(frontend_0_n_55_25), .A1(frontend_0_n_55_7), 
      .A2(frontend_0_n_55_9), .A3(frontend_0_n_55_17), .A4(frontend_0_n_55_24));
  NAND3_X1_LVT frontend_0_i_55_29 (.ZN(frontend_0_n_55_29), .A1(
      frontend_0_n_55_27), .A2(frontend_0_n_55_28), .A3(frontend_0_n_57));
  INV_X1_LVT frontend_0_i_54_0 (.ZN(frontend_0_n_66), .A(
      frontend_0_inst_sext_rdy));
  NAND2_X1_LVT frontend_0_i_55_31 (.ZN(frontend_0_n_55_31), .A1(
      frontend_0_n_55_30), .A2(frontend_0_n_66));
  INV_X1_LVT frontend_0_i_53_1 (.ZN(frontend_0_n_53_0), .A(frontend_0_n_64));
  INV_X1_LVT frontend_0_i_53_2 (.ZN(frontend_0_n_53_1), .A(frontend_0_n_62));
  OAI21_X1_LVT frontend_0_i_53_3 (.ZN(frontend_0_n_65), .A(frontend_0_n_53_0), 
      .B1(frontend_0_n_53_1), .B2(frontend_0_n_63));
  NAND2_X1_LVT frontend_0_i_55_34 (.ZN(frontend_0_n_55_34), .A1(
      frontend_0_n_55_33), .A2(frontend_0_n_65));
  NAND4_X1_LVT frontend_0_i_55_35 (.ZN(frontend_0_e_state_nxt_reg[0]), .A1(
      frontend_0_n_55_25), .A2(frontend_0_n_55_29), .A3(frontend_0_n_55_31), .A4(
      frontend_0_n_55_34));
  DFFS_X1_LVT \frontend_0_e_state_reg[0] (.Q(e_state[0]), .QN(), .CK(cpu_mclk), 
      .D(frontend_0_e_state_nxt_reg[0]), .SN(frontend_0_n_91));
  NAND2_X1_LVT frontend_0_i_32_0 (.ZN(frontend_0_n_32_0), .A1(e_state[0]), .A2(
      e_state[3]));
  NOR3_X1_LVT frontend_0_i_32_1 (.ZN(frontend_0_n_41), .A1(frontend_0_n_32_0), 
      .A2(e_state[1]), .A3(e_state[2]));
  INV_X1_LVT frontend_0_i_33_0 (.ZN(frontend_0_n_33_0), .A(e_state[1]));
  INV_X1_LVT frontend_0_i_33_1 (.ZN(frontend_0_n_33_1), .A(e_state[2]));
  NAND4_X1_LVT frontend_0_i_33_2 (.ZN(frontend_0_n_33_2), .A1(frontend_0_n_33_0), 
      .A2(frontend_0_n_33_1), .A3(e_state[0]), .A4(e_state[3]));
  INV_X1_LVT frontend_0_i_33_3 (.ZN(frontend_0_n_33_3), .A(e_state[0]));
  NAND4_X1_LVT frontend_0_i_33_4 (.ZN(frontend_0_n_33_4), .A1(frontend_0_n_33_3), 
      .A2(frontend_0_n_33_1), .A3(e_state[1]), .A4(e_state[3]));
  NAND2_X1_LVT frontend_0_i_33_5 (.ZN(frontend_0_n_42), .A1(frontend_0_n_33_2), 
      .A2(frontend_0_n_33_4));
  CLKGATETST_X1_LVT frontend_0_clk_gate_exec_dst_wr_reg (.GCK(frontend_0_n_40), 
      .CK(cpu_mclk), .E(frontend_0_n_42), .SE(1'b0));
  DFFR_X1_LVT frontend_0_exec_dst_wr_reg (.Q(frontend_0_exec_dst_wr), .QN(), .CK(
      frontend_0_n_40), .D(frontend_0_n_41), .RN(frontend_0_n_91));
  INV_X1_LVT frontend_0_i_55_42 (.ZN(frontend_0_n_55_41), .A(
      frontend_0_exec_dst_wr));
  NAND2_X1_LVT frontend_0_i_55_56 (.ZN(frontend_0_n_55_54), .A1(
      frontend_0_n_55_41), .A2(frontend_0_exec_jmp));
  INV_X1_LVT frontend_0_i_55_57 (.ZN(frontend_0_n_55_55), .A(frontend_0_n_55_54));
  INV_X1_LVT frontend_0_i_55_58 (.ZN(frontend_0_n_55_56), .A(frontend_0_n_55_16));
  NAND4_X1_LVT frontend_0_i_50_19 (.ZN(frontend_0_n_59), .A1(frontend_0_n_50_16), 
      .A2(frontend_0_n_50_10), .A3(frontend_0_n_50_11), .A4(frontend_0_n_50_13));
  AOI211_X1_LVT frontend_0_i_55_59 (.ZN(frontend_0_n_55_57), .A(
      frontend_0_n_55_55), .B(frontend_0_n_55_56), .C1(frontend_0_n_55_14), .C2(
      frontend_0_n_59));
  NOR2_X1_LVT frontend_0_i_55_60 (.ZN(frontend_0_n_55_58), .A1(
      frontend_0_n_55_57), .A2(frontend_0_n_55_11));
  AND2_X1_LVT frontend_0_i_55_61 (.ZN(frontend_0_n_55_59), .A1(frontend_0_n_55_6), 
      .A2(frontend_0_n_59));
  NOR4_X1_LVT frontend_0_i_55_62 (.ZN(frontend_0_n_55_60), .A1(
      frontend_0_n_55_58), .A2(frontend_0_n_55_59), .A3(frontend_0_n_55_50), .A4(
      frontend_0_n_55_30));
  NOR2_X1_LVT frontend_0_i_55_72 (.ZN(frontend_0_n_55_68), .A1(frontend_0_n_59), 
      .A2(frontend_0_exec_jmp));
  OAI21_X1_LVT frontend_0_i_55_63 (.ZN(frontend_0_e_state_nxt_reg[2]), .A(
      frontend_0_n_55_60), .B1(frontend_0_n_55_26), .B2(frontend_0_n_55_68));
  DFFR_X1_LVT \frontend_0_e_state_reg[2] (.Q(e_state[2]), .QN(), .CK(cpu_mclk), 
      .D(frontend_0_e_state_nxt_reg[2]), .RN(frontend_0_n_91));
  INV_X1_LVT frontend_0_i_55_10 (.ZN(frontend_0_n_55_10), .A(e_state[2]));
  NOR4_X1_LVT frontend_0_i_55_21 (.ZN(frontend_0_n_55_21), .A1(
      frontend_0_n_55_10), .A2(e_state[0]), .A3(e_state[1]), .A4(e_state[3]));
  NOR4_X1_LVT frontend_0_i_55_64 (.ZN(frontend_0_n_55_61), .A1(
      frontend_0_n_55_21), .A2(frontend_0_n_55_36), .A3(frontend_0_n_55_33), .A4(
      frontend_0_n_55_8));
  INV_X1_LVT frontend_0_i_50_20 (.ZN(frontend_0_n_50_17), .A(frontend_0_n_50_6));
  NAND2_X1_LVT frontend_0_i_50_21 (.ZN(frontend_0_n_50_18), .A1(
      frontend_0_n_50_17), .A2(frontend_0_dst_acalc_pre));
  AND4_X1_LVT frontend_0_i_50_22 (.ZN(frontend_0_n_50_19), .A1(frontend_0_n_50_9), 
      .A2(frontend_0_n_50_18), .A3(frontend_0_n_50_11), .A4(frontend_0_n_50_13));
  NAND2_X1_LVT frontend_0_i_50_23 (.ZN(frontend_0_n_60), .A1(frontend_0_n_50_19), 
      .A2(frontend_0_n_50_15));
  INV_X1_LVT frontend_0_i_55_65 (.ZN(frontend_0_n_55_62), .A(frontend_0_n_60));
  NOR2_X1_LVT frontend_0_i_55_66 (.ZN(frontend_0_n_55_63), .A1(
      frontend_0_n_55_62), .A2(frontend_0_exec_jmp));
  OAI21_X1_LVT frontend_0_i_55_67 (.ZN(frontend_0_n_55_64), .A(
      frontend_0_n_55_27), .B1(frontend_0_n_55_63), .B2(frontend_0_exec_jmp));
  OAI211_X1_LVT frontend_0_i_55_68 (.ZN(frontend_0_n_55_65), .A(
      frontend_0_n_55_54), .B(frontend_0_n_55_41), .C1(frontend_0_n_55_42), .C2(
      frontend_0_n_55_62));
  NAND2_X1_LVT frontend_0_i_55_69 (.ZN(frontend_0_n_55_66), .A1(
      frontend_0_n_55_40), .A2(frontend_0_n_55_65));
  NAND2_X1_LVT frontend_0_i_55_70 (.ZN(frontend_0_n_55_67), .A1(
      frontend_0_n_55_6), .A2(frontend_0_n_60));
  NAND4_X1_LVT frontend_0_i_55_71 (.ZN(frontend_0_e_state_nxt_reg[3]), .A1(
      frontend_0_n_55_61), .A2(frontend_0_n_55_64), .A3(frontend_0_n_55_66), .A4(
      frontend_0_n_55_67));
  DFFR_X1_LVT \frontend_0_e_state_reg[3] (.Q(e_state[3]), .QN(), .CK(cpu_mclk), 
      .D(frontend_0_e_state_nxt_reg[3]), .RN(frontend_0_n_91));
  INV_X1_LVT frontend_0_i_58_0 (.ZN(frontend_0_n_58_0), .A(e_state[3]));
  NOR4_X1_LVT frontend_0_i_58_3 (.ZN(frontend_0_n_67), .A1(frontend_0_n_58_0), 
      .A2(frontend_0_n_58_1), .A3(frontend_0_n_58_2), .A4(e_state[1]));
  AND2_X1_LVT frontend_0_i_72_0 (.ZN(frontend_0_n_82), .A1(
      frontend_0_cpu_halt_req), .A2(frontend_0_n_67));
  OAI21_X1_LVT frontend_0_i_72_1 (.ZN(frontend_0_n_72_0), .A(exec_done), .B1(
      frontend_0_cpu_halt_req), .B2(cpuoff));
  INV_X1_LVT frontend_0_i_72_2 (.ZN(frontend_0_n_83), .A(frontend_0_n_72_0));
  NOR2_X1_LVT frontend_0_i_73_0 (.ZN(frontend_0_n_73_0), .A1(frontend_0_n_82), 
      .A2(frontend_0_n_83));
  NOR2_X1_LVT frontend_0_i_73_6 (.ZN(frontend_0_n_86), .A1(frontend_0_n_73_0), 
      .A2(frontend_0_irq_detect));
  NOR3_X1_LVT frontend_0_i_76_13 (.ZN(frontend_0_n_76_12), .A1(frontend_0_n_76_5), 
      .A2(frontend_0_n_76_2), .A3(frontend_0_i_state[2]));
  INV_X1_LVT frontend_0_i_71_0 (.ZN(frontend_0_n_71_0), .A(pc_sw_wr));
  INV_X1_LVT frontend_0_i_64_0 (.ZN(frontend_0_n_64_0), .A(
      frontend_0_dst_acalc_pre));
  NOR2_X1_LVT frontend_0_i_64_1 (.ZN(frontend_0_n_74), .A1(frontend_0_n_64_0), 
      .A2(frontend_0_n_11));
  OR2_X1_LVT frontend_0_i_65_0 (.ZN(frontend_0_n_75), .A1(
      frontend_0_inst_as_nxt[5]), .A2(frontend_0_src_acalc_pre));
  HA_X1_LVT frontend_0_i_66_0 (.CO(frontend_0_inst_sz_nxt[1]), .S(
      frontend_0_inst_sz_nxt[0]), .A(frontend_0_n_74), .B(frontend_0_n_75));
  CLKGATETST_X1_LVT frontend_0_clk_gate_inst_sz_reg (.GCK(frontend_0_n_76), .CK(
      cpu_mclk), .E(frontend_0_decode), .SE(1'b0));
  DFFR_X1_LVT \frontend_0_inst_sz_reg[1] (.Q(frontend_0_inst_sz[1]), .QN(), .CK(
      frontend_0_n_76), .D(frontend_0_inst_sz_nxt[1]), .RN(frontend_0_n_91));
  INV_X1_LVT frontend_0_i_70_0 (.ZN(frontend_0_n_70_0), .A(frontend_0_inst_sz[1]));
  DFFR_X1_LVT \frontend_0_inst_sz_reg[0] (.Q(frontend_0_inst_sz[0]), .QN(), .CK(
      frontend_0_n_76), .D(frontend_0_inst_sz_nxt[0]), .RN(frontend_0_n_91));
  NAND2_X1_LVT frontend_0_i_70_1 (.ZN(frontend_0_n_79), .A1(frontend_0_n_70_0), 
      .A2(frontend_0_inst_sz[0]));
  AND2_X1_LVT frontend_0_i_71_1 (.ZN(frontend_0_n_80), .A1(frontend_0_n_71_0), 
      .A2(frontend_0_n_79));
  AOI221_X1_LVT frontend_0_i_76_16 (.ZN(frontend_0_n_76_14), .A(
      frontend_0_n_76_4), .B1(frontend_0_n_76_6), .B2(frontend_0_n_86), .C1(
      frontend_0_n_76_12), .C2(frontend_0_n_80));
  INV_X1_LVT frontend_0_i_76_17 (.ZN(frontend_0_i_state_nxt_reg[2]), .A(
      frontend_0_n_76_14));
  DFFR_X1_LVT \frontend_0_i_state_reg[2] (.Q(frontend_0_i_state[2]), .QN(), .CK(
      cpu_mclk), .D(frontend_0_i_state_nxt_reg[2]), .RN(frontend_0_n_91));
  OAI33_X1_LVT frontend_0_i_76_9 (.ZN(frontend_0_n_76_8), .A1(frontend_0_n_76_2), 
      .A2(frontend_0_i_state[1]), .A3(frontend_0_i_state[2]), .B1(
      frontend_0_n_76_1), .B2(frontend_0_i_state[0]), .B3(frontend_0_i_state[1]));
  INV_X1_LVT frontend_0_i_76_10 (.ZN(frontend_0_n_76_9), .A(frontend_0_n_76_8));
  INV_X1_LVT frontend_0_i_75_1 (.ZN(frontend_0_n_75_0), .A(frontend_0_n_87));
  NOR2_X1_LVT frontend_0_i_75_2 (.ZN(frontend_0_n_90), .A1(frontend_0_n_75_0), 
      .A2(frontend_0_n_88));
  NAND2_X1_LVT frontend_0_i_76_11 (.ZN(frontend_0_n_76_10), .A1(
      frontend_0_n_76_3), .A2(frontend_0_n_90));
  INV_X1_LVT frontend_0_i_73_1 (.ZN(frontend_0_n_73_1), .A(frontend_0_n_73_0));
  NOR2_X1_LVT frontend_0_i_73_5 (.ZN(frontend_0_n_85), .A1(frontend_0_n_73_1), 
      .A2(frontend_0_irq_detect));
  NAND2_X1_LVT frontend_0_i_76_12 (.ZN(frontend_0_n_76_11), .A1(
      frontend_0_n_76_6), .A2(frontend_0_n_85));
  INV_X1_LVT frontend_0_i_71_2 (.ZN(frontend_0_n_81), .A(frontend_0_n_80));
  NAND2_X1_LVT frontend_0_i_76_14 (.ZN(frontend_0_n_76_13), .A1(
      frontend_0_n_76_12), .A2(frontend_0_n_81));
  NAND4_X1_LVT frontend_0_i_76_15 (.ZN(frontend_0_i_state_nxt_reg[1]), .A1(
      frontend_0_n_76_9), .A2(frontend_0_n_76_10), .A3(frontend_0_n_76_11), .A4(
      frontend_0_n_76_13));
  DFFR_X1_LVT \frontend_0_i_state_reg[1] (.Q(frontend_0_i_state[1]), .QN(), .CK(
      cpu_mclk), .D(frontend_0_i_state_nxt_reg[1]), .RN(frontend_0_n_91));
  NOR3_X1_LVT frontend_0_i_76_0 (.ZN(frontend_0_n_76_0), .A1(
      frontend_0_i_state[0]), .A2(frontend_0_i_state[1]), .A3(
      frontend_0_i_state[2]));
  NOR2_X1_LVT frontend_0_i_68_0 (.ZN(frontend_0_n_77), .A1(exec_done), .A2(
      frontend_0_n_67));
  OR2_X1_LVT frontend_0_i_69_0 (.ZN(frontend_0_n_78), .A1(
      frontend_0_inst_sz_nxt[0]), .A2(frontend_0_inst_sz_nxt[1]));
  INV_X1_LVT frontend_0_i_73_2 (.ZN(frontend_0_n_73_2), .A(frontend_0_n_78));
  OR4_X1_LVT frontend_0_i_73_3 (.ZN(frontend_0_n_73_3), .A1(frontend_0_n_73_1), 
      .A2(frontend_0_n_77), .A3(pc_sw_wr), .A4(frontend_0_n_73_2));
  AOI21_X1_LVT frontend_0_i_73_4 (.ZN(frontend_0_n_84), .A(frontend_0_irq_detect), 
      .B1(frontend_0_n_73_3), .B2(frontend_0_n_73_0));
  AOI211_X1_LVT frontend_0_i_76_7 (.ZN(frontend_0_n_76_7), .A(frontend_0_n_76_0), 
      .B(frontend_0_n_76_4), .C1(frontend_0_n_76_6), .C2(frontend_0_n_84));
  INV_X1_LVT frontend_0_i_76_8 (.ZN(frontend_0_i_state_nxt_reg[0]), .A(
      frontend_0_n_76_7));
  NAND3_X1_LVT frontend_0_i_80_0 (.ZN(frontend_0_n_80_0), .A1(
      frontend_0_i_state_nxt_reg[0]), .A2(frontend_0_i_state_nxt_reg[2]), .A3(
      frontend_0_cpu_halt_req));
  NOR2_X1_LVT frontend_0_i_80_1 (.ZN(frontend_0_n_92), .A1(frontend_0_n_80_0), 
      .A2(frontend_0_i_state_nxt_reg[1]));
  DFFR_X1_LVT frontend_0_cpu_halt_st_reg (.Q(cpu_halt_st), .QN(), .CK(cpu_mclk), 
      .D(frontend_0_n_92), .RN(frontend_0_n_91));
  DFFR_X1_LVT \frontend_0_inst_ad_reg[7] (.Q(inst_ad[7]), .QN(), .CK(
      frontend_0_n_21), .D(1'b0), .RN(frontend_0_n_91));
  DFFR_X1_LVT \frontend_0_inst_ad_reg[5] (.Q(inst_ad[5]), .QN(), .CK(
      frontend_0_n_21), .D(1'b0), .RN(frontend_0_n_91));
  DFFR_X1_LVT \frontend_0_inst_ad_reg[3] (.Q(inst_ad[3]), .QN(), .CK(
      frontend_0_n_21), .D(1'b0), .RN(frontend_0_n_91));
  DFFR_X1_LVT \frontend_0_inst_ad_reg[2] (.Q(inst_ad[2]), .QN(), .CK(
      frontend_0_n_21), .D(1'b0), .RN(frontend_0_n_91));
  DFFR_X1_LVT \frontend_0_inst_ad_reg[0] (.Q(inst_ad[0]), .QN(), .CK(
      frontend_0_n_21), .D(frontend_0_n_18), .RN(frontend_0_n_91));
  INV_X1_LVT frontend_0_i_12_0 (.ZN(frontend_0_n_12_0), .A(
      frontend_0_inst_type_nxt));
  NAND2_X1_LVT frontend_0_i_12_23 (.ZN(frontend_0_n_12_14), .A1(
      frontend_0_n_12_8), .A2(frontend_0_n_12_0));
  NAND3_X1_LVT frontend_0_i_12_5 (.ZN(frontend_0_n_12_5), .A1(frontend_0_n_12_2), 
      .A2(frontend_0_n_12_3), .A3(frontend_0_n_12_4));
  NOR2_X1_LVT frontend_0_i_12_24 (.ZN(frontend_0_inst_as_nxt[9]), .A1(
      frontend_0_n_12_14), .A2(frontend_0_n_12_5));
  NOR2_X1_LVT frontend_0_i_12_25 (.ZN(frontend_0_inst_as_nxt[10]), .A1(
      frontend_0_n_12_14), .A2(frontend_0_n_12_3));
  NOR2_X1_LVT frontend_0_i_12_26 (.ZN(frontend_0_inst_as_nxt[11]), .A1(
      frontend_0_n_12_14), .A2(frontend_0_n_12_2));
  NOR2_X1_LVT frontend_0_i_12_27 (.ZN(frontend_0_inst_as_nxt[12]), .A1(
      frontend_0_n_12_14), .A2(frontend_0_n_12_4));
  NOR4_X1_LVT frontend_0_i_13_0 (.ZN(frontend_0_n_13_0), .A1(
      frontend_0_inst_as_nxt[9]), .A2(frontend_0_inst_as_nxt[10]), .A3(
      frontend_0_inst_as_nxt[11]), .A4(frontend_0_inst_as_nxt[12]));
  NOR3_X1_LVT frontend_0_i_12_21 (.ZN(frontend_0_inst_as_nxt[7]), .A1(
      frontend_0_n_12_13), .A2(frontend_0_n_12_9), .A3(frontend_0_n_12_2));
  NOR3_X1_LVT frontend_0_i_12_22 (.ZN(frontend_0_inst_as_nxt[8]), .A1(
      frontend_0_n_12_13), .A2(frontend_0_n_12_9), .A3(frontend_0_n_12_4));
  NOR2_X1_LVT frontend_0_i_13_1 (.ZN(frontend_0_n_13_1), .A1(
      frontend_0_inst_as_nxt[7]), .A2(frontend_0_inst_as_nxt[8]));
  NAND2_X1_LVT frontend_0_i_13_2 (.ZN(frontend_0_is_const), .A1(
      frontend_0_n_13_0), .A2(frontend_0_n_13_1));
  DFFR_X1_LVT \frontend_0_inst_as_reg[7] (.Q(inst_as[7]), .QN(), .CK(
      frontend_0_n_12), .D(frontend_0_is_const), .RN(frontend_0_n_91));
  DFFR_X1_LVT \frontend_0_inst_as_reg[3] (.Q(inst_as[3]), .QN(), .CK(
      frontend_0_n_12), .D(frontend_0_inst_as_nxt[3]), .RN(frontend_0_n_91));
  DFFR_X1_LVT \frontend_0_inst_as_reg[2] (.Q(inst_as[2]), .QN(), .CK(
      frontend_0_n_12), .D(frontend_0_inst_as_nxt[2]), .RN(frontend_0_n_91));
  OAI21_X1_LVT frontend_0_i_12_10 (.ZN(frontend_0_inst_as_nxt[0]), .A(
      frontend_0_n_12_0), .B1(frontend_0_n_12_5), .B2(frontend_0_n_12_9));
  DFFR_X1_LVT \frontend_0_inst_as_reg[0] (.Q(inst_as[0]), .QN(), .CK(
      frontend_0_n_12), .D(frontend_0_inst_as_nxt[0]), .RN(frontend_0_n_91));
  INV_X1_LVT frontend_0_i_82_1 (.ZN(frontend_0_n_82_1), .A(fe_mdb_in[13]));
  NAND2_X1_LVT frontend_0_i_82_3 (.ZN(frontend_0_n_82_3), .A1(fe_mdb_in[12]), 
      .A2(frontend_0_n_82_1));
  INV_X1_LVT frontend_0_i_82_6 (.ZN(frontend_0_n_82_6), .A(fe_mdb_in[14]));
  NAND2_X1_LVT frontend_0_i_82_9 (.ZN(frontend_0_n_82_9), .A1(frontend_0_n_82_6), 
      .A2(fe_mdb_in[15]));
  NOR2_X1_LVT frontend_0_i_82_16 (.ZN(frontend_0_n_98), .A1(frontend_0_n_82_3), 
      .A2(frontend_0_n_82_9));
  AND2_X1_LVT frontend_0_i_83_5 (.ZN(frontend_0_inst_to_nxt[5]), .A1(
      frontend_0_n_17), .A2(frontend_0_n_98));
  NAND2_X1_LVT frontend_0_i_82_5 (.ZN(frontend_0_n_82_5), .A1(fe_mdb_in[12]), 
      .A2(fe_mdb_in[13]));
  NOR2_X1_LVT frontend_0_i_82_18 (.ZN(frontend_0_n_100), .A1(frontend_0_n_82_5), 
      .A2(frontend_0_n_82_9));
  AND2_X1_LVT frontend_0_i_83_7 (.ZN(frontend_0_inst_to_nxt[7]), .A1(
      frontend_0_n_17), .A2(frontend_0_n_100));
  OR2_X1_LVT frontend_0_i_88_9 (.ZN(frontend_0_inst_alu_nxt[11]), .A1(
      frontend_0_inst_to_nxt[5]), .A2(frontend_0_inst_to_nxt[7]));
  CLKGATETST_X1_LVT frontend_0_clk_gate_inst_alu_reg (.GCK(frontend_0_n_108), 
      .CK(cpu_mclk), .E(frontend_0_decode), .SE(1'b0));
  DFFR_X1_LVT \frontend_0_inst_alu_reg[11] (.Q(inst_alu[11]), .QN(), .CK(
      frontend_0_n_108), .D(frontend_0_inst_alu_nxt[11]), .RN(frontend_0_n_91));
  NOR2_X1_LVT frontend_0_i_25_9 (.ZN(frontend_0_n_24), .A1(frontend_0_n_25_4), 
      .A2(fe_mdb_in[9]));
  AND2_X1_LVT frontend_0_i_26_2 (.ZN(frontend_0_n_32), .A1(frontend_0_n_10), .A2(
      frontend_0_n_24));
  AND2_X1_LVT frontend_0_i_27_3 (.ZN(frontend_0_inst_so_nxt[2]), .A1(
      frontend_0_n_27_0), .A2(frontend_0_n_32));
  NOR2_X1_LVT frontend_0_i_25_7 (.ZN(frontend_0_n_22), .A1(frontend_0_n_25_2), 
      .A2(fe_mdb_in[9]));
  AND2_X1_LVT frontend_0_i_26_0 (.ZN(frontend_0_n_30), .A1(frontend_0_n_22), .A2(
      frontend_0_n_10));
  AND2_X1_LVT frontend_0_i_27_1 (.ZN(frontend_0_inst_so_nxt[0]), .A1(
      frontend_0_n_27_0), .A2(frontend_0_n_30));
  NOR2_X1_LVT frontend_0_i_88_6 (.ZN(frontend_0_n_88_1), .A1(
      frontend_0_inst_so_nxt[2]), .A2(frontend_0_inst_so_nxt[0]));
  INV_X1_LVT frontend_0_i_88_8 (.ZN(frontend_0_inst_alu_nxt[10]), .A(
      frontend_0_n_88_1));
  DFFR_X1_LVT \frontend_0_inst_alu_reg[10] (.Q(inst_alu[10]), .QN(), .CK(
      frontend_0_n_108), .D(frontend_0_inst_alu_nxt[10]), .RN(frontend_0_n_91));
  NAND2_X1_LVT frontend_0_i_82_10 (.ZN(frontend_0_n_82_10), .A1(fe_mdb_in[14]), 
      .A2(fe_mdb_in[15]));
  NOR2_X1_LVT frontend_0_i_82_22 (.ZN(frontend_0_n_104), .A1(frontend_0_n_82_5), 
      .A2(frontend_0_n_82_10));
  AND2_X1_LVT frontend_0_i_83_11 (.ZN(frontend_0_inst_to_nxt[11]), .A1(
      frontend_0_n_17), .A2(frontend_0_n_104));
  OR2_X1_LVT frontend_0_i_87_0 (.ZN(frontend_0_n_107), .A1(
      frontend_0_inst_to_nxt[7]), .A2(frontend_0_inst_to_nxt[11]));
  NOR2_X1_LVT frontend_0_i_25_10 (.ZN(frontend_0_n_25), .A1(frontend_0_n_25_5), 
      .A2(fe_mdb_in[9]));
  AND2_X1_LVT frontend_0_i_26_3 (.ZN(frontend_0_n_33), .A1(frontend_0_n_10), .A2(
      frontend_0_n_25));
  AND2_X1_LVT frontend_0_i_27_4 (.ZN(frontend_0_inst_so_nxt[3]), .A1(
      frontend_0_n_27_0), .A2(frontend_0_n_33));
  OR2_X1_LVT frontend_0_i_88_4 (.ZN(frontend_0_inst_alu_nxt[8]), .A1(
      frontend_0_n_107), .A2(frontend_0_inst_so_nxt[3]));
  INV_X1_LVT frontend_0_i_82_7 (.ZN(frontend_0_n_82_7), .A(fe_mdb_in[15]));
  NAND2_X1_LVT frontend_0_i_82_8 (.ZN(frontend_0_n_82_8), .A1(fe_mdb_in[14]), 
      .A2(frontend_0_n_82_7));
  NOR2_X1_LVT frontend_0_i_82_12 (.ZN(frontend_0_n_94), .A1(frontend_0_n_82_3), 
      .A2(frontend_0_n_82_8));
  AND2_X1_LVT frontend_0_i_83_1 (.ZN(frontend_0_inst_to_nxt[1]), .A1(
      frontend_0_n_17), .A2(frontend_0_n_94));
  INV_X1_LVT frontend_0_i_82_0 (.ZN(frontend_0_n_82_0), .A(fe_mdb_in[12]));
  NAND2_X1_LVT frontend_0_i_82_2 (.ZN(frontend_0_n_82_2), .A1(frontend_0_n_82_0), 
      .A2(frontend_0_n_82_1));
  NOR2_X1_LVT frontend_0_i_82_15 (.ZN(frontend_0_n_97), .A1(frontend_0_n_82_2), 
      .A2(frontend_0_n_82_9));
  AND2_X1_LVT frontend_0_i_83_4 (.ZN(frontend_0_inst_to_nxt[4]), .A1(
      frontend_0_n_17), .A2(frontend_0_n_97));
  OR2_X1_LVT frontend_0_i_84_0 (.ZN(frontend_0_alu_inc), .A1(
      frontend_0_inst_to_nxt[5]), .A2(frontend_0_inst_to_nxt[4]));
  NOR2_X1_LVT frontend_0_i_82_14 (.ZN(frontend_0_n_96), .A1(frontend_0_n_82_5), 
      .A2(frontend_0_n_82_8));
  AND2_X1_LVT frontend_0_i_83_3 (.ZN(frontend_0_inst_to_nxt[3]), .A1(
      frontend_0_n_17), .A2(frontend_0_n_96));
  NAND2_X1_LVT frontend_0_i_82_4 (.ZN(frontend_0_n_82_4), .A1(frontend_0_n_82_0), 
      .A2(fe_mdb_in[13]));
  NOR2_X1_LVT frontend_0_i_82_13 (.ZN(frontend_0_n_95), .A1(frontend_0_n_82_4), 
      .A2(frontend_0_n_82_8));
  AND2_X1_LVT frontend_0_i_83_2 (.ZN(frontend_0_inst_to_nxt[2]), .A1(
      frontend_0_n_17), .A2(frontend_0_n_95));
  OR2_X1_LVT frontend_0_i_85_0 (.ZN(frontend_0_n_105), .A1(
      frontend_0_inst_to_nxt[3]), .A2(frontend_0_inst_to_nxt[2]));
  OR3_X1_LVT frontend_0_i_86_0 (.ZN(frontend_0_n_106), .A1(
      frontend_0_inst_to_nxt[1]), .A2(frontend_0_alu_inc), .A3(frontend_0_n_105));
  NOR2_X1_LVT frontend_0_i_82_21 (.ZN(frontend_0_n_103), .A1(frontend_0_n_82_4), 
      .A2(frontend_0_n_82_10));
  AND2_X1_LVT frontend_0_i_83_10 (.ZN(frontend_0_inst_to_nxt[10]), .A1(
      frontend_0_n_17), .A2(frontend_0_n_103));
  NOR2_X1_LVT frontend_0_i_82_17 (.ZN(frontend_0_n_99), .A1(frontend_0_n_82_4), 
      .A2(frontend_0_n_82_9));
  AND2_X1_LVT frontend_0_i_83_6 (.ZN(frontend_0_inst_to_nxt[6]), .A1(
      frontend_0_n_17), .A2(frontend_0_n_99));
  NOR4_X1_LVT frontend_0_i_88_5 (.ZN(frontend_0_n_88_0), .A1(
      frontend_0_inst_alu_nxt[8]), .A2(frontend_0_n_106), .A3(
      frontend_0_inst_to_nxt[10]), .A4(frontend_0_inst_to_nxt[6]));
  NAND2_X1_LVT frontend_0_i_88_7 (.ZN(frontend_0_inst_alu_nxt[9]), .A1(
      frontend_0_n_88_0), .A2(frontend_0_n_88_1));
  DFFR_X1_LVT \frontend_0_inst_alu_reg[9] (.Q(inst_alu[9]), .QN(), .CK(
      frontend_0_n_108), .D(frontend_0_inst_alu_nxt[9]), .RN(frontend_0_n_91));
  DFFR_X1_LVT \frontend_0_inst_alu_reg[8] (.Q(inst_alu[8]), .QN(), .CK(
      frontend_0_n_108), .D(frontend_0_inst_alu_nxt[8]), .RN(frontend_0_n_91));
  DFFR_X1_LVT \frontend_0_inst_alu_reg[7] (.Q(inst_alu[7]), .QN(), .CK(
      frontend_0_n_108), .D(frontend_0_inst_to_nxt[6]), .RN(frontend_0_n_91));
  DFFR_X1_LVT \frontend_0_inst_alu_reg[6] (.Q(inst_alu[6]), .QN(), .CK(
      frontend_0_n_108), .D(frontend_0_inst_to_nxt[10]), .RN(frontend_0_n_91));
  NOR2_X1_LVT frontend_0_i_82_20 (.ZN(frontend_0_n_102), .A1(frontend_0_n_82_3), 
      .A2(frontend_0_n_82_10));
  AND2_X1_LVT frontend_0_i_83_9 (.ZN(frontend_0_inst_to_nxt[9]), .A1(
      frontend_0_n_17), .A2(frontend_0_n_102));
  DFFR_X1_LVT \frontend_0_inst_alu_reg[5] (.Q(inst_alu[5]), .QN(), .CK(
      frontend_0_n_108), .D(frontend_0_inst_to_nxt[9]), .RN(frontend_0_n_91));
  NOR2_X1_LVT frontend_0_i_82_19 (.ZN(frontend_0_n_101), .A1(frontend_0_n_82_2), 
      .A2(frontend_0_n_82_10));
  AND2_X1_LVT frontend_0_i_83_8 (.ZN(frontend_0_inst_to_nxt[8]), .A1(
      frontend_0_n_17), .A2(frontend_0_n_101));
  OR2_X1_LVT frontend_0_i_88_3 (.ZN(frontend_0_inst_alu_nxt[4]), .A1(
      frontend_0_inst_to_nxt[8]), .A2(frontend_0_n_107));
  DFFR_X1_LVT \frontend_0_inst_alu_reg[4] (.Q(inst_alu[4]), .QN(), .CK(
      frontend_0_n_108), .D(frontend_0_inst_alu_nxt[4]), .RN(frontend_0_n_91));
  OR2_X1_LVT frontend_0_i_88_2 (.ZN(frontend_0_inst_alu_nxt[3]), .A1(
      frontend_0_n_49), .A2(frontend_0_n_106));
  DFFR_X1_LVT \frontend_0_inst_alu_reg[3] (.Q(inst_alu[3]), .QN(), .CK(
      frontend_0_n_108), .D(frontend_0_inst_alu_nxt[3]), .RN(frontend_0_n_91));
  OR2_X1_LVT frontend_0_i_88_1 (.ZN(frontend_0_inst_alu_nxt[2]), .A1(
      frontend_0_inst_to_nxt[6]), .A2(frontend_0_n_105));
  DFFR_X1_LVT \frontend_0_inst_alu_reg[2] (.Q(inst_alu[2]), .QN(), .CK(
      frontend_0_n_108), .D(frontend_0_inst_alu_nxt[2]), .RN(frontend_0_n_91));
  DFFR_X1_LVT \frontend_0_inst_alu_reg[1] (.Q(inst_alu[1]), .QN(), .CK(
      frontend_0_n_108), .D(frontend_0_alu_inc), .RN(frontend_0_n_91));
  OR3_X1_LVT frontend_0_i_88_0 (.ZN(frontend_0_inst_alu_nxt[0]), .A1(
      frontend_0_inst_to_nxt[3]), .A2(frontend_0_alu_inc), .A3(
      frontend_0_inst_to_nxt[8]));
  DFFR_X1_LVT \frontend_0_inst_alu_reg[0] (.Q(inst_alu[0]), .QN(), .CK(
      frontend_0_n_108), .D(frontend_0_inst_alu_nxt[0]), .RN(frontend_0_n_91));
  NAND3_X1_LVT frontend_0_i_91_0 (.ZN(frontend_0_n_91_0), .A1(fe_mdb_in[6]), .A2(
      frontend_0_n_0), .A3(frontend_0_n_9));
  NOR2_X1_LVT frontend_0_i_91_1 (.ZN(frontend_0_n_110), .A1(frontend_0_n_91_0), 
      .A2(frontend_0_inst_type_nxt));
  CLKGATETST_X1_LVT frontend_0_clk_gate_inst_bw_reg (.GCK(frontend_0_n_109), .CK(
      cpu_mclk), .E(frontend_0_decode), .SE(1'b0));
  DFFR_X1_LVT frontend_0_inst_bw_reg (.Q(inst_bw), .QN(), .CK(frontend_0_n_109), 
      .D(frontend_0_n_110), .RN(frontend_0_n_91));
  DFFR_X1_LVT \frontend_0_inst_type_reg[1] (.Q(inst_type[1]), .QN(), .CK(
      frontend_0_n_43), .D(frontend_0_inst_type_nxt), .RN(frontend_0_n_91));
  NOR2_X1_LVT frontend_0_i_97_0 (.ZN(frontend_0_n_97_0), .A1(inst_type[1]), .A2(
      cpu_halt_st));
  INV_X1_LVT frontend_0_i_97_1 (.ZN(frontend_0_n_97_1), .A(frontend_0_n_97_0));
  DFFR_X1_LVT \frontend_0_inst_so_reg[7] (.Q(inst_so[7]), .QN(), .CK(
      frontend_0_n_38), .D(frontend_0_inst_so_nxt[7]), .RN(frontend_0_n_91));
  OR2_X1_LVT frontend_0_i_96_0 (.ZN(frontend_0_n_144), .A1(inst_so[7]), .A2(
      frontend_0_n_39));
  NOR2_X1_LVT frontend_0_i_97_2 (.ZN(frontend_0_n_97_2), .A1(frontend_0_n_97_1), 
      .A2(frontend_0_n_144));
  CLKGATETST_X1_LVT frontend_0_clk_gate_inst_dest_bin_reg (.GCK(frontend_0_n_111), 
      .CK(cpu_mclk), .E(frontend_0_decode), .SE(1'b0));
  DFFR_X1_LVT \frontend_0_inst_dest_bin_reg[0] (.Q(frontend_0_inst_dest_bin[0]), 
      .QN(), .CK(frontend_0_n_111), .D(fe_mdb_in[0]), .RN(frontend_0_n_91));
  DFFR_X1_LVT \frontend_0_inst_dest_bin_reg[1] (.Q(frontend_0_inst_dest_bin[1]), 
      .QN(), .CK(frontend_0_n_111), .D(fe_mdb_in[1]), .RN(frontend_0_n_91));
  NAND2_X1_LVT frontend_0_i_94_5 (.ZN(frontend_0_n_94_5), .A1(
      frontend_0_inst_dest_bin[0]), .A2(frontend_0_inst_dest_bin[1]));
  DFFR_X1_LVT \frontend_0_inst_dest_bin_reg[2] (.Q(frontend_0_inst_dest_bin[2]), 
      .QN(), .CK(frontend_0_n_111), .D(fe_mdb_in[2]), .RN(frontend_0_n_91));
  DFFR_X1_LVT \frontend_0_inst_dest_bin_reg[3] (.Q(frontend_0_inst_dest_bin[3]), 
      .QN(), .CK(frontend_0_n_111), .D(fe_mdb_in[3]), .RN(frontend_0_n_91));
  NAND2_X1_LVT frontend_0_i_94_11 (.ZN(frontend_0_n_94_11), .A1(
      frontend_0_inst_dest_bin[2]), .A2(frontend_0_inst_dest_bin[3]));
  NOR2_X1_LVT frontend_0_i_94_27 (.ZN(frontend_0_n_127), .A1(frontend_0_n_94_5), 
      .A2(frontend_0_n_94_11));
  NAND2_X1_LVT frontend_0_i_95_5 (.ZN(frontend_0_n_95_5), .A1(dbg_mem_addr[0]), 
      .A2(dbg_mem_addr[1]));
  NAND2_X1_LVT frontend_0_i_95_11 (.ZN(frontend_0_n_95_11), .A1(dbg_mem_addr[2]), 
      .A2(dbg_mem_addr[3]));
  NOR2_X1_LVT frontend_0_i_95_27 (.ZN(frontend_0_n_143), .A1(frontend_0_n_95_5), 
      .A2(frontend_0_n_95_11));
  AOI22_X1_LVT frontend_0_i_97_34 (.ZN(frontend_0_n_97_19), .A1(
      frontend_0_n_97_2), .A2(frontend_0_n_127), .B1(cpu_halt_st), .B2(
      frontend_0_n_143));
  INV_X1_LVT frontend_0_i_97_35 (.ZN(inst_dest[15]), .A(frontend_0_n_97_19));
  INV_X1_LVT frontend_0_i_94_0 (.ZN(frontend_0_n_94_0), .A(
      frontend_0_inst_dest_bin[0]));
  NAND2_X1_LVT frontend_0_i_94_4 (.ZN(frontend_0_n_94_4), .A1(frontend_0_n_94_0), 
      .A2(frontend_0_inst_dest_bin[1]));
  NOR2_X1_LVT frontend_0_i_94_26 (.ZN(frontend_0_n_126), .A1(frontend_0_n_94_4), 
      .A2(frontend_0_n_94_11));
  INV_X1_LVT frontend_0_i_95_0 (.ZN(frontend_0_n_95_0), .A(dbg_mem_addr[0]));
  NAND2_X1_LVT frontend_0_i_95_4 (.ZN(frontend_0_n_95_4), .A1(frontend_0_n_95_0), 
      .A2(dbg_mem_addr[1]));
  NOR2_X1_LVT frontend_0_i_95_26 (.ZN(frontend_0_n_142), .A1(frontend_0_n_95_4), 
      .A2(frontend_0_n_95_11));
  AOI22_X1_LVT frontend_0_i_97_32 (.ZN(frontend_0_n_97_18), .A1(
      frontend_0_n_97_2), .A2(frontend_0_n_126), .B1(cpu_halt_st), .B2(
      frontend_0_n_142));
  INV_X1_LVT frontend_0_i_97_33 (.ZN(inst_dest[14]), .A(frontend_0_n_97_18));
  INV_X1_LVT frontend_0_i_94_1 (.ZN(frontend_0_n_94_1), .A(
      frontend_0_inst_dest_bin[1]));
  NAND2_X1_LVT frontend_0_i_94_3 (.ZN(frontend_0_n_94_3), .A1(
      frontend_0_inst_dest_bin[0]), .A2(frontend_0_n_94_1));
  NOR2_X1_LVT frontend_0_i_94_25 (.ZN(frontend_0_n_125), .A1(frontend_0_n_94_3), 
      .A2(frontend_0_n_94_11));
  INV_X1_LVT frontend_0_i_95_1 (.ZN(frontend_0_n_95_1), .A(dbg_mem_addr[1]));
  NAND2_X1_LVT frontend_0_i_95_3 (.ZN(frontend_0_n_95_3), .A1(dbg_mem_addr[0]), 
      .A2(frontend_0_n_95_1));
  NOR2_X1_LVT frontend_0_i_95_25 (.ZN(frontend_0_n_141), .A1(frontend_0_n_95_3), 
      .A2(frontend_0_n_95_11));
  AOI22_X1_LVT frontend_0_i_97_30 (.ZN(frontend_0_n_97_17), .A1(
      frontend_0_n_97_2), .A2(frontend_0_n_125), .B1(cpu_halt_st), .B2(
      frontend_0_n_141));
  INV_X1_LVT frontend_0_i_97_31 (.ZN(inst_dest[13]), .A(frontend_0_n_97_17));
  NAND2_X1_LVT frontend_0_i_94_2 (.ZN(frontend_0_n_94_2), .A1(frontend_0_n_94_0), 
      .A2(frontend_0_n_94_1));
  NOR2_X1_LVT frontend_0_i_94_24 (.ZN(frontend_0_n_124), .A1(frontend_0_n_94_2), 
      .A2(frontend_0_n_94_11));
  NAND2_X1_LVT frontend_0_i_95_2 (.ZN(frontend_0_n_95_2), .A1(frontend_0_n_95_0), 
      .A2(frontend_0_n_95_1));
  NOR2_X1_LVT frontend_0_i_95_24 (.ZN(frontend_0_n_140), .A1(frontend_0_n_95_2), 
      .A2(frontend_0_n_95_11));
  AOI22_X1_LVT frontend_0_i_97_28 (.ZN(frontend_0_n_97_16), .A1(
      frontend_0_n_97_2), .A2(frontend_0_n_124), .B1(cpu_halt_st), .B2(
      frontend_0_n_140));
  INV_X1_LVT frontend_0_i_97_29 (.ZN(inst_dest[12]), .A(frontend_0_n_97_16));
  INV_X1_LVT frontend_0_i_94_6 (.ZN(frontend_0_n_94_6), .A(
      frontend_0_inst_dest_bin[2]));
  NAND2_X1_LVT frontend_0_i_94_10 (.ZN(frontend_0_n_94_10), .A1(
      frontend_0_n_94_6), .A2(frontend_0_inst_dest_bin[3]));
  NOR2_X1_LVT frontend_0_i_94_23 (.ZN(frontend_0_n_123), .A1(frontend_0_n_94_5), 
      .A2(frontend_0_n_94_10));
  INV_X1_LVT frontend_0_i_95_6 (.ZN(frontend_0_n_95_6), .A(dbg_mem_addr[2]));
  NAND2_X1_LVT frontend_0_i_95_10 (.ZN(frontend_0_n_95_10), .A1(
      frontend_0_n_95_6), .A2(dbg_mem_addr[3]));
  NOR2_X1_LVT frontend_0_i_95_23 (.ZN(frontend_0_n_139), .A1(frontend_0_n_95_5), 
      .A2(frontend_0_n_95_10));
  AOI22_X1_LVT frontend_0_i_97_26 (.ZN(frontend_0_n_97_15), .A1(
      frontend_0_n_97_2), .A2(frontend_0_n_123), .B1(cpu_halt_st), .B2(
      frontend_0_n_139));
  INV_X1_LVT frontend_0_i_97_27 (.ZN(inst_dest[11]), .A(frontend_0_n_97_15));
  NOR2_X1_LVT frontend_0_i_94_22 (.ZN(frontend_0_n_122), .A1(frontend_0_n_94_4), 
      .A2(frontend_0_n_94_10));
  NOR2_X1_LVT frontend_0_i_95_22 (.ZN(frontend_0_n_138), .A1(frontend_0_n_95_4), 
      .A2(frontend_0_n_95_10));
  AOI22_X1_LVT frontend_0_i_97_24 (.ZN(frontend_0_n_97_14), .A1(
      frontend_0_n_97_2), .A2(frontend_0_n_122), .B1(cpu_halt_st), .B2(
      frontend_0_n_138));
  INV_X1_LVT frontend_0_i_97_25 (.ZN(inst_dest[10]), .A(frontend_0_n_97_14));
  NOR2_X1_LVT frontend_0_i_94_21 (.ZN(frontend_0_n_121), .A1(frontend_0_n_94_3), 
      .A2(frontend_0_n_94_10));
  NOR2_X1_LVT frontend_0_i_95_21 (.ZN(frontend_0_n_137), .A1(frontend_0_n_95_3), 
      .A2(frontend_0_n_95_10));
  AOI22_X1_LVT frontend_0_i_97_22 (.ZN(frontend_0_n_97_13), .A1(
      frontend_0_n_97_2), .A2(frontend_0_n_121), .B1(cpu_halt_st), .B2(
      frontend_0_n_137));
  INV_X1_LVT frontend_0_i_97_23 (.ZN(inst_dest[9]), .A(frontend_0_n_97_13));
  NOR2_X1_LVT frontend_0_i_94_20 (.ZN(frontend_0_n_120), .A1(frontend_0_n_94_2), 
      .A2(frontend_0_n_94_10));
  NOR2_X1_LVT frontend_0_i_95_20 (.ZN(frontend_0_n_136), .A1(frontend_0_n_95_2), 
      .A2(frontend_0_n_95_10));
  AOI22_X1_LVT frontend_0_i_97_20 (.ZN(frontend_0_n_97_12), .A1(
      frontend_0_n_97_2), .A2(frontend_0_n_120), .B1(cpu_halt_st), .B2(
      frontend_0_n_136));
  INV_X1_LVT frontend_0_i_97_21 (.ZN(inst_dest[8]), .A(frontend_0_n_97_12));
  INV_X1_LVT frontend_0_i_94_7 (.ZN(frontend_0_n_94_7), .A(
      frontend_0_inst_dest_bin[3]));
  NAND2_X1_LVT frontend_0_i_94_9 (.ZN(frontend_0_n_94_9), .A1(
      frontend_0_inst_dest_bin[2]), .A2(frontend_0_n_94_7));
  NOR2_X1_LVT frontend_0_i_94_19 (.ZN(frontend_0_n_119), .A1(frontend_0_n_94_5), 
      .A2(frontend_0_n_94_9));
  INV_X1_LVT frontend_0_i_95_7 (.ZN(frontend_0_n_95_7), .A(dbg_mem_addr[3]));
  NAND2_X1_LVT frontend_0_i_95_9 (.ZN(frontend_0_n_95_9), .A1(dbg_mem_addr[2]), 
      .A2(frontend_0_n_95_7));
  NOR2_X1_LVT frontend_0_i_95_19 (.ZN(frontend_0_n_135), .A1(frontend_0_n_95_5), 
      .A2(frontend_0_n_95_9));
  AOI22_X1_LVT frontend_0_i_97_18 (.ZN(frontend_0_n_97_11), .A1(
      frontend_0_n_97_2), .A2(frontend_0_n_119), .B1(cpu_halt_st), .B2(
      frontend_0_n_135));
  INV_X1_LVT frontend_0_i_97_19 (.ZN(inst_dest[7]), .A(frontend_0_n_97_11));
  NOR2_X1_LVT frontend_0_i_94_18 (.ZN(frontend_0_n_118), .A1(frontend_0_n_94_4), 
      .A2(frontend_0_n_94_9));
  NOR2_X1_LVT frontend_0_i_95_18 (.ZN(frontend_0_n_134), .A1(frontend_0_n_95_4), 
      .A2(frontend_0_n_95_9));
  AOI22_X1_LVT frontend_0_i_97_16 (.ZN(frontend_0_n_97_10), .A1(
      frontend_0_n_97_2), .A2(frontend_0_n_118), .B1(cpu_halt_st), .B2(
      frontend_0_n_134));
  INV_X1_LVT frontend_0_i_97_17 (.ZN(inst_dest[6]), .A(frontend_0_n_97_10));
  NOR2_X1_LVT frontend_0_i_94_17 (.ZN(frontend_0_n_117), .A1(frontend_0_n_94_3), 
      .A2(frontend_0_n_94_9));
  NOR2_X1_LVT frontend_0_i_95_17 (.ZN(frontend_0_n_133), .A1(frontend_0_n_95_3), 
      .A2(frontend_0_n_95_9));
  AOI22_X1_LVT frontend_0_i_97_14 (.ZN(frontend_0_n_97_9), .A1(frontend_0_n_97_2), 
      .A2(frontend_0_n_117), .B1(cpu_halt_st), .B2(frontend_0_n_133));
  INV_X1_LVT frontend_0_i_97_15 (.ZN(inst_dest[5]), .A(frontend_0_n_97_9));
  NOR2_X1_LVT frontend_0_i_94_16 (.ZN(frontend_0_n_116), .A1(frontend_0_n_94_2), 
      .A2(frontend_0_n_94_9));
  NOR2_X1_LVT frontend_0_i_95_16 (.ZN(frontend_0_n_132), .A1(frontend_0_n_95_2), 
      .A2(frontend_0_n_95_9));
  AOI22_X1_LVT frontend_0_i_97_12 (.ZN(frontend_0_n_97_8), .A1(frontend_0_n_97_2), 
      .A2(frontend_0_n_116), .B1(cpu_halt_st), .B2(frontend_0_n_132));
  INV_X1_LVT frontend_0_i_97_13 (.ZN(inst_dest[4]), .A(frontend_0_n_97_8));
  NAND2_X1_LVT frontend_0_i_94_8 (.ZN(frontend_0_n_94_8), .A1(frontend_0_n_94_6), 
      .A2(frontend_0_n_94_7));
  NOR2_X1_LVT frontend_0_i_94_15 (.ZN(frontend_0_n_115), .A1(frontend_0_n_94_5), 
      .A2(frontend_0_n_94_8));
  NAND2_X1_LVT frontend_0_i_95_8 (.ZN(frontend_0_n_95_8), .A1(frontend_0_n_95_6), 
      .A2(frontend_0_n_95_7));
  NOR2_X1_LVT frontend_0_i_95_15 (.ZN(frontend_0_n_131), .A1(frontend_0_n_95_5), 
      .A2(frontend_0_n_95_8));
  AOI22_X1_LVT frontend_0_i_97_10 (.ZN(frontend_0_n_97_7), .A1(frontend_0_n_97_2), 
      .A2(frontend_0_n_115), .B1(cpu_halt_st), .B2(frontend_0_n_131));
  INV_X1_LVT frontend_0_i_97_11 (.ZN(inst_dest[3]), .A(frontend_0_n_97_7));
  NOR2_X1_LVT frontend_0_i_94_14 (.ZN(frontend_0_n_114), .A1(frontend_0_n_94_4), 
      .A2(frontend_0_n_94_8));
  NOR2_X1_LVT frontend_0_i_95_14 (.ZN(frontend_0_n_130), .A1(frontend_0_n_95_4), 
      .A2(frontend_0_n_95_8));
  AOI22_X1_LVT frontend_0_i_97_8 (.ZN(frontend_0_n_97_6), .A1(frontend_0_n_97_2), 
      .A2(frontend_0_n_114), .B1(cpu_halt_st), .B2(frontend_0_n_130));
  INV_X1_LVT frontend_0_i_97_9 (.ZN(inst_dest[2]), .A(frontend_0_n_97_6));
  NOR2_X1_LVT frontend_0_i_94_13 (.ZN(frontend_0_n_113), .A1(frontend_0_n_94_3), 
      .A2(frontend_0_n_94_8));
  NOR2_X1_LVT frontend_0_i_95_13 (.ZN(frontend_0_n_129), .A1(frontend_0_n_95_3), 
      .A2(frontend_0_n_95_8));
  AOI222_X1_LVT frontend_0_i_97_6 (.ZN(frontend_0_n_97_5), .A1(frontend_0_n_97_2), 
      .A2(frontend_0_n_113), .B1(frontend_0_n_97_0), .B2(frontend_0_n_144), .C1(
      cpu_halt_st), .C2(frontend_0_n_129));
  INV_X1_LVT frontend_0_i_97_7 (.ZN(inst_dest[1]), .A(frontend_0_n_97_5));
  NOR2_X1_LVT frontend_0_i_94_12 (.ZN(frontend_0_n_112), .A1(frontend_0_n_94_2), 
      .A2(frontend_0_n_94_8));
  INV_X1_LVT frontend_0_i_97_3 (.ZN(frontend_0_n_97_3), .A(cpu_halt_st));
  NOR2_X1_LVT frontend_0_i_95_12 (.ZN(frontend_0_n_128), .A1(frontend_0_n_95_2), 
      .A2(frontend_0_n_95_8));
  AOI222_X1_LVT frontend_0_i_97_4 (.ZN(frontend_0_n_97_4), .A1(frontend_0_n_97_2), 
      .A2(frontend_0_n_112), .B1(frontend_0_n_97_3), .B2(inst_type[1]), .C1(
      frontend_0_n_128), .C2(cpu_halt_st));
  INV_X1_LVT frontend_0_i_97_5 (.ZN(inst_dest[0]), .A(frontend_0_n_97_4));
  INV_X1_LVT frontend_0_i_99_6 (.ZN(frontend_0_n_99_4), .A(fe_mdb_in[3]));
  XNOR2_X1_LVT frontend_0_i_99_19 (.ZN(frontend_0_n_99_17), .A(fe_mdb_in[15]), 
      .B(frontend_0_n_99_4));
  INV_X1_LVT frontend_0_i_98_0 (.ZN(frontend_0_n_98_0), .A(
      frontend_0_i_state_nxt_reg[2]));
  OR3_X1_LVT frontend_0_i_98_1 (.ZN(frontend_0_n_98_1), .A1(frontend_0_n_98_0), 
      .A2(frontend_0_i_state_nxt_reg[0]), .A3(frontend_0_i_state_nxt_reg[1]));
  INV_X1_LVT frontend_0_i_98_2 (.ZN(frontend_0_n_98_2), .A(inst_as[4]));
  AND4_X1_LVT frontend_0_i_98_3 (.ZN(frontend_0_n_98_3), .A1(frontend_0_n_98_1), 
      .A2(frontend_0_n_98_2), .A3(frontend_0_n_6), .A4(inst_ad[4]));
  AOI221_X1_LVT frontend_0_i_98_4 (.ZN(frontend_0_n_98_4), .A(frontend_0_n_98_3), 
      .B1(frontend_0_n_6), .B2(inst_as[4]), .C1(frontend_0_n_7), .C2(inst_ad[4]));
  INV_X1_LVT frontend_0_i_98_5 (.ZN(frontend_0_n_145), .A(frontend_0_n_98_4));
  INV_X1_LVT frontend_0_i_99_3 (.ZN(frontend_0_n_99_2), .A(fe_mdb_in[1]));
  NAND2_X1_LVT frontend_0_i_99_2 (.ZN(frontend_0_n_99_1), .A1(frontend_0_n_145), 
      .A2(frontend_0_n_99_2));
  OR2_X1_LVT frontend_0_i_99_5 (.ZN(frontend_0_n_99_3), .A1(fe_mdb_in[2]), .A2(
      frontend_0_n_99_1));
  HA_X1_LVT frontend_0_i_99_7 (.CO(frontend_0_n_99_5), .S(frontend_0_ext_nxt[3]), 
      .A(frontend_0_n_99_4), .B(frontend_0_n_99_3));
  FA_X1_LVT frontend_0_i_99_8 (.CO(frontend_0_n_99_6), .S(frontend_0_ext_nxt[4]), 
      .A(fe_mdb_in[4]), .B(frontend_0_n_99_4), .CI(frontend_0_n_99_5));
  FA_X1_LVT frontend_0_i_99_9 (.CO(frontend_0_n_99_7), .S(frontend_0_ext_nxt[5]), 
      .A(fe_mdb_in[5]), .B(frontend_0_n_99_4), .CI(frontend_0_n_99_6));
  FA_X1_LVT frontend_0_i_99_10 (.CO(frontend_0_n_99_8), .S(frontend_0_ext_nxt[6]), 
      .A(fe_mdb_in[6]), .B(frontend_0_n_99_4), .CI(frontend_0_n_99_7));
  FA_X1_LVT frontend_0_i_99_11 (.CO(frontend_0_n_99_9), .S(frontend_0_ext_nxt[7]), 
      .A(fe_mdb_in[7]), .B(frontend_0_n_99_4), .CI(frontend_0_n_99_8));
  FA_X1_LVT frontend_0_i_99_12 (.CO(frontend_0_n_99_10), .S(
      frontend_0_ext_nxt[8]), .A(fe_mdb_in[8]), .B(frontend_0_n_99_4), .CI(
      frontend_0_n_99_9));
  FA_X1_LVT frontend_0_i_99_13 (.CO(frontend_0_n_99_11), .S(
      frontend_0_ext_nxt[9]), .A(fe_mdb_in[9]), .B(frontend_0_n_99_4), .CI(
      frontend_0_n_99_10));
  FA_X1_LVT frontend_0_i_99_14 (.CO(frontend_0_n_99_12), .S(
      frontend_0_ext_nxt[10]), .A(fe_mdb_in[10]), .B(frontend_0_n_99_4), .CI(
      frontend_0_n_99_11));
  FA_X1_LVT frontend_0_i_99_15 (.CO(frontend_0_n_99_13), .S(
      frontend_0_ext_nxt[11]), .A(fe_mdb_in[11]), .B(frontend_0_n_99_4), .CI(
      frontend_0_n_99_12));
  FA_X1_LVT frontend_0_i_99_16 (.CO(frontend_0_n_99_14), .S(
      frontend_0_ext_nxt[12]), .A(fe_mdb_in[12]), .B(frontend_0_n_99_4), .CI(
      frontend_0_n_99_13));
  FA_X1_LVT frontend_0_i_99_17 (.CO(frontend_0_n_99_15), .S(
      frontend_0_ext_nxt[13]), .A(fe_mdb_in[13]), .B(frontend_0_n_99_4), .CI(
      frontend_0_n_99_14));
  FA_X1_LVT frontend_0_i_99_18 (.CO(frontend_0_n_99_16), .S(
      frontend_0_ext_nxt[14]), .A(fe_mdb_in[14]), .B(frontend_0_n_99_4), .CI(
      frontend_0_n_99_15));
  XNOR2_X1_LVT frontend_0_i_99_20 (.ZN(frontend_0_ext_nxt[15]), .A(
      frontend_0_n_99_17), .B(frontend_0_n_99_16));
  INV_X1_LVT frontend_0_i_101_0 (.ZN(frontend_0_n_101_0), .A(
      frontend_0_i_state[2]));
  NOR3_X1_LVT frontend_0_i_101_1 (.ZN(frontend_0_n_101_1), .A1(
      frontend_0_n_101_0), .A2(frontend_0_i_state[0]), .A3(frontend_0_i_state[1]));
  OR2_X1_LVT frontend_0_i_101_2 (.ZN(frontend_0_n_147), .A1(frontend_0_n_101_1), 
      .A2(frontend_0_n_13));
  CLKGATETST_X1_LVT frontend_0_clk_gate_inst_dext_reg (.GCK(frontend_0_n_146), 
      .CK(cpu_mclk), .E(frontend_0_n_147), .SE(1'b0));
  DFFR_X1_LVT \frontend_0_inst_dext_reg[15] (.Q(inst_dext[15]), .QN(), .CK(
      frontend_0_n_146), .D(frontend_0_ext_nxt[15]), .RN(frontend_0_n_91));
  DFFR_X1_LVT \frontend_0_inst_dext_reg[14] (.Q(inst_dext[14]), .QN(), .CK(
      frontend_0_n_146), .D(frontend_0_ext_nxt[14]), .RN(frontend_0_n_91));
  DFFR_X1_LVT \frontend_0_inst_dext_reg[13] (.Q(inst_dext[13]), .QN(), .CK(
      frontend_0_n_146), .D(frontend_0_ext_nxt[13]), .RN(frontend_0_n_91));
  DFFR_X1_LVT \frontend_0_inst_dext_reg[12] (.Q(inst_dext[12]), .QN(), .CK(
      frontend_0_n_146), .D(frontend_0_ext_nxt[12]), .RN(frontend_0_n_91));
  DFFR_X1_LVT \frontend_0_inst_dext_reg[11] (.Q(inst_dext[11]), .QN(), .CK(
      frontend_0_n_146), .D(frontend_0_ext_nxt[11]), .RN(frontend_0_n_91));
  DFFR_X1_LVT \frontend_0_inst_dext_reg[10] (.Q(inst_dext[10]), .QN(), .CK(
      frontend_0_n_146), .D(frontend_0_ext_nxt[10]), .RN(frontend_0_n_91));
  DFFR_X1_LVT \frontend_0_inst_dext_reg[9] (.Q(inst_dext[9]), .QN(), .CK(
      frontend_0_n_146), .D(frontend_0_ext_nxt[9]), .RN(frontend_0_n_91));
  DFFR_X1_LVT \frontend_0_inst_dext_reg[8] (.Q(inst_dext[8]), .QN(), .CK(
      frontend_0_n_146), .D(frontend_0_ext_nxt[8]), .RN(frontend_0_n_91));
  DFFR_X1_LVT \frontend_0_inst_dext_reg[7] (.Q(inst_dext[7]), .QN(), .CK(
      frontend_0_n_146), .D(frontend_0_ext_nxt[7]), .RN(frontend_0_n_91));
  DFFR_X1_LVT \frontend_0_inst_dext_reg[6] (.Q(inst_dext[6]), .QN(), .CK(
      frontend_0_n_146), .D(frontend_0_ext_nxt[6]), .RN(frontend_0_n_91));
  DFFR_X1_LVT \frontend_0_inst_dext_reg[5] (.Q(inst_dext[5]), .QN(), .CK(
      frontend_0_n_146), .D(frontend_0_ext_nxt[5]), .RN(frontend_0_n_91));
  DFFR_X1_LVT \frontend_0_inst_dext_reg[4] (.Q(inst_dext[4]), .QN(), .CK(
      frontend_0_n_146), .D(frontend_0_ext_nxt[4]), .RN(frontend_0_n_91));
  DFFR_X1_LVT \frontend_0_inst_dext_reg[3] (.Q(inst_dext[3]), .QN(), .CK(
      frontend_0_n_146), .D(frontend_0_ext_nxt[3]), .RN(frontend_0_n_91));
  XNOR2_X1_LVT frontend_0_i_99_4 (.ZN(frontend_0_ext_nxt[2]), .A(fe_mdb_in[2]), 
      .B(frontend_0_n_99_1));
  DFFR_X1_LVT \frontend_0_inst_dext_reg[2] (.Q(inst_dext[2]), .QN(), .CK(
      frontend_0_n_146), .D(frontend_0_ext_nxt[2]), .RN(frontend_0_n_91));
  XNOR2_X1_LVT frontend_0_i_99_0 (.ZN(frontend_0_n_99_0), .A(frontend_0_n_145), 
      .B(fe_mdb_in[1]));
  INV_X1_LVT frontend_0_i_99_1 (.ZN(frontend_0_ext_nxt[1]), .A(frontend_0_n_99_0));
  DFFR_X1_LVT \frontend_0_inst_dext_reg[1] (.Q(inst_dext[1]), .QN(), .CK(
      frontend_0_n_146), .D(frontend_0_ext_nxt[1]), .RN(frontend_0_n_91));
  DFFR_X1_LVT \frontend_0_inst_dext_reg[0] (.Q(inst_dext[0]), .QN(), .CK(
      frontend_0_n_146), .D(fe_mdb_in[0]), .RN(frontend_0_n_91));
  CLKGATETST_X1_LVT frontend_0_clk_gate_inst_irq_rst_reg (.GCK(frontend_0_n_148), 
      .CK(cpu_mclk), .E(exec_done), .SE(1'b0));
  DFFS_X1_LVT frontend_0_inst_irq_rst_reg (.Q(inst_irq_rst), .QN(), .CK(
      frontend_0_n_148), .D(1'b0), .SN(frontend_0_n_91));
  CLKGATETST_X1_LVT frontend_0_clk_gate_inst_jmp_bin_reg (.GCK(frontend_0_n_149), 
      .CK(cpu_mclk), .E(frontend_0_decode), .SE(1'b0));
  DFFR_X1_LVT \frontend_0_inst_jmp_bin_reg[0] (.Q(frontend_0_inst_jmp_bin[0]), 
      .QN(), .CK(frontend_0_n_149), .D(fe_mdb_in[10]), .RN(frontend_0_n_91));
  DFFR_X1_LVT \frontend_0_inst_jmp_bin_reg[1] (.Q(frontend_0_inst_jmp_bin[1]), 
      .QN(), .CK(frontend_0_n_149), .D(fe_mdb_in[11]), .RN(frontend_0_n_91));
  NAND2_X1_LVT frontend_0_i_105_5 (.ZN(frontend_0_n_105_5), .A1(
      frontend_0_inst_jmp_bin[0]), .A2(frontend_0_inst_jmp_bin[1]));
  DFFR_X1_LVT \frontend_0_inst_jmp_bin_reg[2] (.Q(frontend_0_inst_jmp_bin[2]), 
      .QN(), .CK(frontend_0_n_149), .D(fe_mdb_in[12]), .RN(frontend_0_n_91));
  INV_X1_LVT frontend_0_i_105_6 (.ZN(frontend_0_n_105_6), .A(
      frontend_0_inst_jmp_bin[2]));
  NOR2_X1_LVT frontend_0_i_105_14 (.ZN(frontend_0_n_157), .A1(frontend_0_n_105_5), 
      .A2(frontend_0_n_105_6));
  AND2_X1_LVT frontend_0_i_106_7 (.ZN(inst_jmp[7]), .A1(inst_type[1]), .A2(
      frontend_0_n_157));
  INV_X1_LVT frontend_0_i_105_0 (.ZN(frontend_0_n_105_0), .A(
      frontend_0_inst_jmp_bin[0]));
  NAND2_X1_LVT frontend_0_i_105_4 (.ZN(frontend_0_n_105_4), .A1(
      frontend_0_n_105_0), .A2(frontend_0_inst_jmp_bin[1]));
  NOR2_X1_LVT frontend_0_i_105_13 (.ZN(frontend_0_n_156), .A1(frontend_0_n_105_4), 
      .A2(frontend_0_n_105_6));
  AND2_X1_LVT frontend_0_i_106_6 (.ZN(inst_jmp[6]), .A1(inst_type[1]), .A2(
      frontend_0_n_156));
  INV_X1_LVT frontend_0_i_105_1 (.ZN(frontend_0_n_105_1), .A(
      frontend_0_inst_jmp_bin[1]));
  NAND2_X1_LVT frontend_0_i_105_3 (.ZN(frontend_0_n_105_3), .A1(
      frontend_0_inst_jmp_bin[0]), .A2(frontend_0_n_105_1));
  NOR2_X1_LVT frontend_0_i_105_12 (.ZN(frontend_0_n_155), .A1(frontend_0_n_105_3), 
      .A2(frontend_0_n_105_6));
  AND2_X1_LVT frontend_0_i_106_5 (.ZN(inst_jmp[5]), .A1(inst_type[1]), .A2(
      frontend_0_n_155));
  NAND2_X1_LVT frontend_0_i_105_2 (.ZN(frontend_0_n_105_2), .A1(
      frontend_0_n_105_0), .A2(frontend_0_n_105_1));
  NOR2_X1_LVT frontend_0_i_105_11 (.ZN(frontend_0_n_154), .A1(frontend_0_n_105_2), 
      .A2(frontend_0_n_105_6));
  AND2_X1_LVT frontend_0_i_106_4 (.ZN(inst_jmp[4]), .A1(inst_type[1]), .A2(
      frontend_0_n_154));
  NOR2_X1_LVT frontend_0_i_105_10 (.ZN(frontend_0_n_153), .A1(frontend_0_n_105_5), 
      .A2(frontend_0_inst_jmp_bin[2]));
  AND2_X1_LVT frontend_0_i_106_3 (.ZN(inst_jmp[3]), .A1(inst_type[1]), .A2(
      frontend_0_n_153));
  NOR2_X1_LVT frontend_0_i_105_9 (.ZN(frontend_0_n_152), .A1(frontend_0_n_105_4), 
      .A2(frontend_0_inst_jmp_bin[2]));
  AND2_X1_LVT frontend_0_i_106_2 (.ZN(inst_jmp[2]), .A1(inst_type[1]), .A2(
      frontend_0_n_152));
  NOR2_X1_LVT frontend_0_i_105_8 (.ZN(frontend_0_n_151), .A1(frontend_0_n_105_3), 
      .A2(frontend_0_inst_jmp_bin[2]));
  AND2_X1_LVT frontend_0_i_106_1 (.ZN(inst_jmp[1]), .A1(inst_type[1]), .A2(
      frontend_0_n_151));
  NOR2_X1_LVT frontend_0_i_105_7 (.ZN(frontend_0_n_150), .A1(frontend_0_n_105_2), 
      .A2(frontend_0_inst_jmp_bin[2]));
  AND2_X1_LVT frontend_0_i_106_0 (.ZN(inst_jmp[0]), .A1(frontend_0_n_150), .A2(
      inst_type[1]));
  NOR2_X1_LVT frontend_0_i_82_11 (.ZN(frontend_0_n_93), .A1(frontend_0_n_82_2), 
      .A2(frontend_0_n_82_8));
  AND2_X1_LVT frontend_0_i_83_0 (.ZN(frontend_0_inst_to_nxt[0]), .A1(
      frontend_0_n_17), .A2(frontend_0_n_93));
  CLKGATETST_X1_LVT frontend_0_clk_gate_inst_mov_reg (.GCK(frontend_0_n_158), 
      .CK(cpu_mclk), .E(frontend_0_decode), .SE(1'b0));
  DFFR_X1_LVT frontend_0_inst_mov_reg (.Q(inst_mov), .QN(), .CK(frontend_0_n_158), 
      .D(frontend_0_inst_to_nxt[0]), .RN(frontend_0_n_91));
  AND2_X1_LVT frontend_0_i_110_33 (.ZN(frontend_0_n_110_23), .A1(
      frontend_0_inst_type_nxt), .A2(fe_mdb_in[9]));
  AND2_X1_LVT frontend_0_i_110_14 (.ZN(frontend_0_n_110_10), .A1(
      frontend_0_is_const), .A2(frontend_0_inst_as_nxt[12]));
  NOR2_X1_LVT frontend_0_i_110_0 (.ZN(frontend_0_n_110_0), .A1(
      frontend_0_inst_type_nxt), .A2(frontend_0_is_const));
  AOI211_X1_LVT frontend_0_i_110_49 (.ZN(frontend_0_n_110_34), .A(
      frontend_0_n_110_23), .B(frontend_0_n_110_10), .C1(frontend_0_n_110_0), 
      .C2(frontend_0_ext_nxt[15]));
  INV_X1_LVT frontend_0_i_110_2 (.ZN(frontend_0_n_110_2), .A(frontend_0_decode));
  INV_X1_LVT frontend_0_i_110_50 (.ZN(frontend_0_n_110_35), .A(
      frontend_0_ext_nxt[15]));
  OAI22_X1_LVT frontend_0_i_110_51 (.ZN(frontend_0_n_179), .A1(
      frontend_0_n_110_34), .A2(frontend_0_n_110_2), .B1(frontend_0_decode), .B2(
      frontend_0_n_110_35));
  NOR2_X1_LVT frontend_0_i_111_0 (.ZN(frontend_0_n_111_0), .A1(
      frontend_0_inst_type_nxt), .A2(frontend_0_is_const));
  INV_X1_LVT frontend_0_i_111_4 (.ZN(frontend_0_n_111_3), .A(frontend_0_n_111_0));
  NOR2_X1_LVT frontend_0_i_111_5 (.ZN(frontend_0_n_111_4), .A1(
      frontend_0_inst_sext_rdy), .A2(frontend_0_n_111_3));
  INV_X1_LVT frontend_0_i_111_1 (.ZN(frontend_0_n_111_1), .A(frontend_0_decode));
  INV_X1_LVT frontend_0_i_111_2 (.ZN(frontend_0_n_111_2), .A(
      frontend_0_inst_sext_rdy));
  OAI22_X1_LVT frontend_0_i_111_3 (.ZN(frontend_0_n_180), .A1(frontend_0_n_111_4), 
      .A2(frontend_0_n_111_1), .B1(frontend_0_decode), .B2(frontend_0_n_111_2));
  CLKGATETST_X1_LVT frontend_0_clk_gate_inst_sext_reg (.GCK(frontend_0_n_163), 
      .CK(cpu_mclk), .E(frontend_0_n_180), .SE(1'b0));
  DFFR_X1_LVT \frontend_0_inst_sext_reg[15] (.Q(inst_sext[15]), .QN(), .CK(
      frontend_0_n_163), .D(frontend_0_n_179), .RN(frontend_0_n_91));
  AOI211_X1_LVT frontend_0_i_110_46 (.ZN(frontend_0_n_110_32), .A(
      frontend_0_n_110_23), .B(frontend_0_n_110_10), .C1(frontend_0_n_110_0), 
      .C2(frontend_0_ext_nxt[14]));
  INV_X1_LVT frontend_0_i_110_47 (.ZN(frontend_0_n_110_33), .A(
      frontend_0_ext_nxt[14]));
  OAI22_X1_LVT frontend_0_i_110_48 (.ZN(frontend_0_n_178), .A1(
      frontend_0_n_110_32), .A2(frontend_0_n_110_2), .B1(frontend_0_decode), .B2(
      frontend_0_n_110_33));
  DFFR_X1_LVT \frontend_0_inst_sext_reg[14] (.Q(inst_sext[14]), .QN(), .CK(
      frontend_0_n_163), .D(frontend_0_n_178), .RN(frontend_0_n_91));
  AOI211_X1_LVT frontend_0_i_110_43 (.ZN(frontend_0_n_110_30), .A(
      frontend_0_n_110_23), .B(frontend_0_n_110_10), .C1(frontend_0_n_110_0), 
      .C2(frontend_0_ext_nxt[13]));
  INV_X1_LVT frontend_0_i_110_44 (.ZN(frontend_0_n_110_31), .A(
      frontend_0_ext_nxt[13]));
  OAI22_X1_LVT frontend_0_i_110_45 (.ZN(frontend_0_n_177), .A1(
      frontend_0_n_110_30), .A2(frontend_0_n_110_2), .B1(frontend_0_decode), .B2(
      frontend_0_n_110_31));
  DFFR_X1_LVT \frontend_0_inst_sext_reg[13] (.Q(inst_sext[13]), .QN(), .CK(
      frontend_0_n_163), .D(frontend_0_n_177), .RN(frontend_0_n_91));
  AOI211_X1_LVT frontend_0_i_110_40 (.ZN(frontend_0_n_110_28), .A(
      frontend_0_n_110_23), .B(frontend_0_n_110_10), .C1(frontend_0_n_110_0), 
      .C2(frontend_0_ext_nxt[12]));
  INV_X1_LVT frontend_0_i_110_41 (.ZN(frontend_0_n_110_29), .A(
      frontend_0_ext_nxt[12]));
  OAI22_X1_LVT frontend_0_i_110_42 (.ZN(frontend_0_n_176), .A1(
      frontend_0_n_110_28), .A2(frontend_0_n_110_2), .B1(frontend_0_decode), .B2(
      frontend_0_n_110_29));
  DFFR_X1_LVT \frontend_0_inst_sext_reg[12] (.Q(inst_sext[12]), .QN(), .CK(
      frontend_0_n_163), .D(frontend_0_n_176), .RN(frontend_0_n_91));
  AOI211_X1_LVT frontend_0_i_110_37 (.ZN(frontend_0_n_110_26), .A(
      frontend_0_n_110_23), .B(frontend_0_n_110_10), .C1(frontend_0_n_110_0), 
      .C2(frontend_0_ext_nxt[11]));
  INV_X1_LVT frontend_0_i_110_38 (.ZN(frontend_0_n_110_27), .A(
      frontend_0_ext_nxt[11]));
  OAI22_X1_LVT frontend_0_i_110_39 (.ZN(frontend_0_n_175), .A1(
      frontend_0_n_110_26), .A2(frontend_0_n_110_2), .B1(frontend_0_decode), .B2(
      frontend_0_n_110_27));
  DFFR_X1_LVT \frontend_0_inst_sext_reg[11] (.Q(inst_sext[11]), .QN(), .CK(
      frontend_0_n_163), .D(frontend_0_n_175), .RN(frontend_0_n_91));
  AOI211_X1_LVT frontend_0_i_110_34 (.ZN(frontend_0_n_110_24), .A(
      frontend_0_n_110_23), .B(frontend_0_n_110_10), .C1(frontend_0_n_110_0), 
      .C2(frontend_0_ext_nxt[10]));
  INV_X1_LVT frontend_0_i_110_35 (.ZN(frontend_0_n_110_25), .A(
      frontend_0_ext_nxt[10]));
  OAI22_X1_LVT frontend_0_i_110_36 (.ZN(frontend_0_n_174), .A1(
      frontend_0_n_110_24), .A2(frontend_0_n_110_2), .B1(frontend_0_decode), .B2(
      frontend_0_n_110_25));
  DFFR_X1_LVT \frontend_0_inst_sext_reg[10] (.Q(inst_sext[10]), .QN(), .CK(
      frontend_0_n_163), .D(frontend_0_n_174), .RN(frontend_0_n_91));
  AOI221_X1_LVT frontend_0_i_110_30 (.ZN(frontend_0_n_110_21), .A(
      frontend_0_n_110_10), .B1(frontend_0_inst_type_nxt), .B2(fe_mdb_in[8]), 
      .C1(frontend_0_n_110_0), .C2(frontend_0_ext_nxt[9]));
  INV_X1_LVT frontend_0_i_110_31 (.ZN(frontend_0_n_110_22), .A(
      frontend_0_ext_nxt[9]));
  OAI22_X1_LVT frontend_0_i_110_32 (.ZN(frontend_0_n_173), .A1(
      frontend_0_n_110_21), .A2(frontend_0_n_110_2), .B1(frontend_0_decode), .B2(
      frontend_0_n_110_22));
  DFFR_X1_LVT \frontend_0_inst_sext_reg[9] (.Q(inst_sext[9]), .QN(), .CK(
      frontend_0_n_163), .D(frontend_0_n_173), .RN(frontend_0_n_91));
  AOI221_X1_LVT frontend_0_i_110_27 (.ZN(frontend_0_n_110_19), .A(
      frontend_0_n_110_10), .B1(frontend_0_inst_type_nxt), .B2(fe_mdb_in[7]), 
      .C1(frontend_0_n_110_0), .C2(frontend_0_ext_nxt[8]));
  INV_X1_LVT frontend_0_i_110_28 (.ZN(frontend_0_n_110_20), .A(
      frontend_0_ext_nxt[8]));
  OAI22_X1_LVT frontend_0_i_110_29 (.ZN(frontend_0_n_172), .A1(
      frontend_0_n_110_19), .A2(frontend_0_n_110_2), .B1(frontend_0_decode), .B2(
      frontend_0_n_110_20));
  DFFR_X1_LVT \frontend_0_inst_sext_reg[8] (.Q(inst_sext[8]), .QN(), .CK(
      frontend_0_n_163), .D(frontend_0_n_172), .RN(frontend_0_n_91));
  AOI221_X1_LVT frontend_0_i_110_24 (.ZN(frontend_0_n_110_17), .A(
      frontend_0_n_110_10), .B1(frontend_0_inst_type_nxt), .B2(fe_mdb_in[6]), 
      .C1(frontend_0_n_110_0), .C2(frontend_0_ext_nxt[7]));
  INV_X1_LVT frontend_0_i_110_25 (.ZN(frontend_0_n_110_18), .A(
      frontend_0_ext_nxt[7]));
  OAI22_X1_LVT frontend_0_i_110_26 (.ZN(frontend_0_n_171), .A1(
      frontend_0_n_110_17), .A2(frontend_0_n_110_2), .B1(frontend_0_decode), .B2(
      frontend_0_n_110_18));
  DFFR_X1_LVT \frontend_0_inst_sext_reg[7] (.Q(inst_sext[7]), .QN(), .CK(
      frontend_0_n_163), .D(frontend_0_n_171), .RN(frontend_0_n_91));
  AOI221_X1_LVT frontend_0_i_110_21 (.ZN(frontend_0_n_110_15), .A(
      frontend_0_n_110_10), .B1(frontend_0_inst_type_nxt), .B2(fe_mdb_in[5]), 
      .C1(frontend_0_n_110_0), .C2(frontend_0_ext_nxt[6]));
  INV_X1_LVT frontend_0_i_110_22 (.ZN(frontend_0_n_110_16), .A(
      frontend_0_ext_nxt[6]));
  OAI22_X1_LVT frontend_0_i_110_23 (.ZN(frontend_0_n_170), .A1(
      frontend_0_n_110_15), .A2(frontend_0_n_110_2), .B1(frontend_0_decode), .B2(
      frontend_0_n_110_16));
  DFFR_X1_LVT \frontend_0_inst_sext_reg[6] (.Q(inst_sext[6]), .QN(), .CK(
      frontend_0_n_163), .D(frontend_0_n_170), .RN(frontend_0_n_91));
  AOI221_X1_LVT frontend_0_i_110_18 (.ZN(frontend_0_n_110_13), .A(
      frontend_0_n_110_10), .B1(frontend_0_inst_type_nxt), .B2(fe_mdb_in[4]), 
      .C1(frontend_0_n_110_0), .C2(frontend_0_ext_nxt[5]));
  INV_X1_LVT frontend_0_i_110_19 (.ZN(frontend_0_n_110_14), .A(
      frontend_0_ext_nxt[5]));
  OAI22_X1_LVT frontend_0_i_110_20 (.ZN(frontend_0_n_169), .A1(
      frontend_0_n_110_13), .A2(frontend_0_n_110_2), .B1(frontend_0_decode), .B2(
      frontend_0_n_110_14));
  DFFR_X1_LVT \frontend_0_inst_sext_reg[5] (.Q(inst_sext[5]), .QN(), .CK(
      frontend_0_n_163), .D(frontend_0_n_169), .RN(frontend_0_n_91));
  AOI221_X1_LVT frontend_0_i_110_15 (.ZN(frontend_0_n_110_11), .A(
      frontend_0_n_110_10), .B1(frontend_0_inst_type_nxt), .B2(fe_mdb_in[3]), 
      .C1(frontend_0_n_110_0), .C2(frontend_0_ext_nxt[4]));
  INV_X1_LVT frontend_0_i_110_16 (.ZN(frontend_0_n_110_12), .A(
      frontend_0_ext_nxt[4]));
  OAI22_X1_LVT frontend_0_i_110_17 (.ZN(frontend_0_n_168), .A1(
      frontend_0_n_110_11), .A2(frontend_0_n_110_2), .B1(frontend_0_decode), .B2(
      frontend_0_n_110_12));
  DFFR_X1_LVT \frontend_0_inst_sext_reg[4] (.Q(inst_sext[4]), .QN(), .CK(
      frontend_0_n_163), .D(frontend_0_n_168), .RN(frontend_0_n_91));
  OR2_X1_LVT frontend_0_i_108_3 (.ZN(frontend_0_n_162), .A1(
      frontend_0_inst_as_nxt[12]), .A2(frontend_0_inst_as_nxt[8]));
  AOI222_X1_LVT frontend_0_i_110_11 (.ZN(frontend_0_n_110_8), .A1(
      frontend_0_n_110_0), .A2(frontend_0_ext_nxt[3]), .B1(frontend_0_is_const), 
      .B2(frontend_0_n_162), .C1(frontend_0_inst_type_nxt), .C2(fe_mdb_in[2]));
  INV_X1_LVT frontend_0_i_110_12 (.ZN(frontend_0_n_110_9), .A(
      frontend_0_ext_nxt[3]));
  OAI22_X1_LVT frontend_0_i_110_13 (.ZN(frontend_0_n_167), .A1(
      frontend_0_n_110_8), .A2(frontend_0_n_110_2), .B1(frontend_0_decode), .B2(
      frontend_0_n_110_9));
  DFFR_X1_LVT \frontend_0_inst_sext_reg[3] (.Q(inst_sext[3]), .QN(), .CK(
      frontend_0_n_163), .D(frontend_0_n_167), .RN(frontend_0_n_91));
  OR2_X1_LVT frontend_0_i_108_2 (.ZN(frontend_0_n_161), .A1(
      frontend_0_inst_as_nxt[12]), .A2(frontend_0_inst_as_nxt[7]));
  AOI222_X1_LVT frontend_0_i_110_8 (.ZN(frontend_0_n_110_6), .A1(
      frontend_0_n_110_0), .A2(frontend_0_ext_nxt[2]), .B1(frontend_0_is_const), 
      .B2(frontend_0_n_161), .C1(frontend_0_inst_type_nxt), .C2(fe_mdb_in[1]));
  INV_X1_LVT frontend_0_i_110_9 (.ZN(frontend_0_n_110_7), .A(
      frontend_0_ext_nxt[2]));
  OAI22_X1_LVT frontend_0_i_110_10 (.ZN(frontend_0_n_166), .A1(
      frontend_0_n_110_6), .A2(frontend_0_n_110_2), .B1(frontend_0_decode), .B2(
      frontend_0_n_110_7));
  DFFR_X1_LVT \frontend_0_inst_sext_reg[2] (.Q(inst_sext[2]), .QN(), .CK(
      frontend_0_n_163), .D(frontend_0_n_166), .RN(frontend_0_n_91));
  OR2_X1_LVT frontend_0_i_108_1 (.ZN(frontend_0_n_160), .A1(
      frontend_0_inst_as_nxt[12]), .A2(frontend_0_inst_as_nxt[11]));
  AOI222_X1_LVT frontend_0_i_110_5 (.ZN(frontend_0_n_110_4), .A1(
      frontend_0_n_110_0), .A2(frontend_0_ext_nxt[1]), .B1(frontend_0_is_const), 
      .B2(frontend_0_n_160), .C1(frontend_0_inst_type_nxt), .C2(fe_mdb_in[0]));
  INV_X1_LVT frontend_0_i_110_6 (.ZN(frontend_0_n_110_5), .A(
      frontend_0_ext_nxt[1]));
  OAI22_X1_LVT frontend_0_i_110_7 (.ZN(frontend_0_n_165), .A1(frontend_0_n_110_4), 
      .A2(frontend_0_n_110_2), .B1(frontend_0_decode), .B2(frontend_0_n_110_5));
  DFFR_X1_LVT \frontend_0_inst_sext_reg[1] (.Q(inst_sext[1]), .QN(), .CK(
      frontend_0_n_163), .D(frontend_0_n_165), .RN(frontend_0_n_91));
  OR2_X1_LVT frontend_0_i_108_0 (.ZN(frontend_0_n_159), .A1(
      frontend_0_inst_as_nxt[12]), .A2(frontend_0_inst_as_nxt[10]));
  AOI22_X1_LVT frontend_0_i_110_1 (.ZN(frontend_0_n_110_1), .A1(
      frontend_0_n_110_0), .A2(fe_mdb_in[0]), .B1(frontend_0_n_159), .B2(
      frontend_0_is_const));
  INV_X1_LVT frontend_0_i_110_3 (.ZN(frontend_0_n_110_3), .A(fe_mdb_in[0]));
  OAI22_X1_LVT frontend_0_i_110_4 (.ZN(frontend_0_n_164), .A1(frontend_0_n_110_1), 
      .A2(frontend_0_n_110_2), .B1(frontend_0_decode), .B2(frontend_0_n_110_3));
  DFFR_X1_LVT \frontend_0_inst_sext_reg[0] (.Q(inst_sext[0]), .QN(), .CK(
      frontend_0_n_163), .D(frontend_0_n_164), .RN(frontend_0_n_91));
  DFFR_X1_LVT \frontend_0_inst_so_reg[3] (.Q(inst_so[3]), .QN(), .CK(
      frontend_0_n_38), .D(frontend_0_inst_so_nxt[3]), .RN(frontend_0_n_91));
  DFFR_X1_LVT \frontend_0_inst_so_reg[2] (.Q(inst_so[2]), .QN(), .CK(
      frontend_0_n_38), .D(frontend_0_inst_so_nxt[2]), .RN(frontend_0_n_91));
  NOR2_X1_LVT frontend_0_i_25_8 (.ZN(frontend_0_n_23), .A1(frontend_0_n_25_3), 
      .A2(fe_mdb_in[9]));
  AND2_X1_LVT frontend_0_i_26_1 (.ZN(frontend_0_n_31), .A1(frontend_0_n_10), .A2(
      frontend_0_n_23));
  AND2_X1_LVT frontend_0_i_27_2 (.ZN(frontend_0_inst_so_nxt[1]), .A1(
      frontend_0_n_27_0), .A2(frontend_0_n_31));
  DFFR_X1_LVT \frontend_0_inst_so_reg[1] (.Q(inst_so[1]), .QN(), .CK(
      frontend_0_n_38), .D(frontend_0_inst_so_nxt[1]), .RN(frontend_0_n_91));
  DFFR_X1_LVT \frontend_0_inst_so_reg[0] (.Q(inst_so[0]), .QN(), .CK(
      frontend_0_n_38), .D(frontend_0_inst_so_nxt[0]), .RN(frontend_0_n_91));
  DFFR_X1_LVT \frontend_0_inst_type_reg[2] (.Q(inst_type[2]), .QN(), .CK(
      frontend_0_n_43), .D(frontend_0_n_17), .RN(frontend_0_n_91));
  NOR2_X1_LVT frontend_0_i_115_0 (.ZN(frontend_0_n_115_0), .A1(inst_so[6]), .A2(
      inst_type[2]));
  INV_X1_LVT frontend_0_i_115_1 (.ZN(frontend_0_n_115_1), .A(inst_so[7]));
  AND3_X1_LVT frontend_0_i_115_2 (.ZN(frontend_0_n_115_2), .A1(
      frontend_0_n_115_0), .A2(frontend_0_n_115_1), .A3(inst_type[0]));
  CLKGATETST_X1_LVT frontend_0_clk_gate_inst_src_bin_reg (.GCK(frontend_0_n_181), 
      .CK(cpu_mclk), .E(frontend_0_decode), .SE(1'b0));
  DFFR_X1_LVT \frontend_0_inst_src_bin_reg[0] (.Q(frontend_0_inst_src_bin[0]), 
      .QN(), .CK(frontend_0_n_181), .D(fe_mdb_in[8]), .RN(frontend_0_n_91));
  DFFR_X1_LVT \frontend_0_inst_src_bin_reg[1] (.Q(frontend_0_inst_src_bin[1]), 
      .QN(), .CK(frontend_0_n_181), .D(fe_mdb_in[9]), .RN(frontend_0_n_91));
  NAND2_X1_LVT frontend_0_i_114_5 (.ZN(frontend_0_n_114_5), .A1(
      frontend_0_inst_src_bin[0]), .A2(frontend_0_inst_src_bin[1]));
  DFFR_X1_LVT \frontend_0_inst_src_bin_reg[2] (.Q(frontend_0_inst_src_bin[2]), 
      .QN(), .CK(frontend_0_n_181), .D(fe_mdb_in[10]), .RN(frontend_0_n_91));
  DFFR_X1_LVT \frontend_0_inst_src_bin_reg[3] (.Q(frontend_0_inst_src_bin[3]), 
      .QN(), .CK(frontend_0_n_181), .D(fe_mdb_in[11]), .RN(frontend_0_n_91));
  NAND2_X1_LVT frontend_0_i_114_11 (.ZN(frontend_0_n_114_11), .A1(
      frontend_0_inst_src_bin[2]), .A2(frontend_0_inst_src_bin[3]));
  NOR2_X1_LVT frontend_0_i_114_27 (.ZN(frontend_0_n_197), .A1(frontend_0_n_114_5), 
      .A2(frontend_0_n_114_11));
  AOI22_X1_LVT frontend_0_i_115_34 (.ZN(frontend_0_n_115_19), .A1(
      frontend_0_n_115_2), .A2(frontend_0_n_127), .B1(inst_type[2]), .B2(
      frontend_0_n_197));
  INV_X1_LVT frontend_0_i_115_35 (.ZN(inst_src[15]), .A(frontend_0_n_115_19));
  INV_X1_LVT frontend_0_i_114_0 (.ZN(frontend_0_n_114_0), .A(
      frontend_0_inst_src_bin[0]));
  NAND2_X1_LVT frontend_0_i_114_4 (.ZN(frontend_0_n_114_4), .A1(
      frontend_0_n_114_0), .A2(frontend_0_inst_src_bin[1]));
  NOR2_X1_LVT frontend_0_i_114_26 (.ZN(frontend_0_n_196), .A1(frontend_0_n_114_4), 
      .A2(frontend_0_n_114_11));
  AOI22_X1_LVT frontend_0_i_115_32 (.ZN(frontend_0_n_115_18), .A1(
      frontend_0_n_115_2), .A2(frontend_0_n_126), .B1(inst_type[2]), .B2(
      frontend_0_n_196));
  INV_X1_LVT frontend_0_i_115_33 (.ZN(inst_src[14]), .A(frontend_0_n_115_18));
  INV_X1_LVT frontend_0_i_114_1 (.ZN(frontend_0_n_114_1), .A(
      frontend_0_inst_src_bin[1]));
  NAND2_X1_LVT frontend_0_i_114_3 (.ZN(frontend_0_n_114_3), .A1(
      frontend_0_inst_src_bin[0]), .A2(frontend_0_n_114_1));
  NOR2_X1_LVT frontend_0_i_114_25 (.ZN(frontend_0_n_195), .A1(frontend_0_n_114_3), 
      .A2(frontend_0_n_114_11));
  AOI22_X1_LVT frontend_0_i_115_30 (.ZN(frontend_0_n_115_17), .A1(
      frontend_0_n_115_2), .A2(frontend_0_n_125), .B1(inst_type[2]), .B2(
      frontend_0_n_195));
  INV_X1_LVT frontend_0_i_115_31 (.ZN(inst_src[13]), .A(frontend_0_n_115_17));
  NAND2_X1_LVT frontend_0_i_114_2 (.ZN(frontend_0_n_114_2), .A1(
      frontend_0_n_114_0), .A2(frontend_0_n_114_1));
  NOR2_X1_LVT frontend_0_i_114_24 (.ZN(frontend_0_n_194), .A1(frontend_0_n_114_2), 
      .A2(frontend_0_n_114_11));
  AOI22_X1_LVT frontend_0_i_115_28 (.ZN(frontend_0_n_115_16), .A1(
      frontend_0_n_115_2), .A2(frontend_0_n_124), .B1(inst_type[2]), .B2(
      frontend_0_n_194));
  INV_X1_LVT frontend_0_i_115_29 (.ZN(inst_src[12]), .A(frontend_0_n_115_16));
  INV_X1_LVT frontend_0_i_114_6 (.ZN(frontend_0_n_114_6), .A(
      frontend_0_inst_src_bin[2]));
  NAND2_X1_LVT frontend_0_i_114_10 (.ZN(frontend_0_n_114_10), .A1(
      frontend_0_n_114_6), .A2(frontend_0_inst_src_bin[3]));
  NOR2_X1_LVT frontend_0_i_114_23 (.ZN(frontend_0_n_193), .A1(frontend_0_n_114_5), 
      .A2(frontend_0_n_114_10));
  AOI22_X1_LVT frontend_0_i_115_26 (.ZN(frontend_0_n_115_15), .A1(
      frontend_0_n_115_2), .A2(frontend_0_n_123), .B1(inst_type[2]), .B2(
      frontend_0_n_193));
  INV_X1_LVT frontend_0_i_115_27 (.ZN(inst_src[11]), .A(frontend_0_n_115_15));
  NOR2_X1_LVT frontend_0_i_114_22 (.ZN(frontend_0_n_192), .A1(frontend_0_n_114_4), 
      .A2(frontend_0_n_114_10));
  AOI22_X1_LVT frontend_0_i_115_24 (.ZN(frontend_0_n_115_14), .A1(
      frontend_0_n_115_2), .A2(frontend_0_n_122), .B1(inst_type[2]), .B2(
      frontend_0_n_192));
  INV_X1_LVT frontend_0_i_115_25 (.ZN(inst_src[10]), .A(frontend_0_n_115_14));
  NOR2_X1_LVT frontend_0_i_114_21 (.ZN(frontend_0_n_191), .A1(frontend_0_n_114_3), 
      .A2(frontend_0_n_114_10));
  AOI22_X1_LVT frontend_0_i_115_22 (.ZN(frontend_0_n_115_13), .A1(
      frontend_0_n_115_2), .A2(frontend_0_n_121), .B1(inst_type[2]), .B2(
      frontend_0_n_191));
  INV_X1_LVT frontend_0_i_115_23 (.ZN(inst_src[9]), .A(frontend_0_n_115_13));
  NOR2_X1_LVT frontend_0_i_114_20 (.ZN(frontend_0_n_190), .A1(frontend_0_n_114_2), 
      .A2(frontend_0_n_114_10));
  AOI22_X1_LVT frontend_0_i_115_20 (.ZN(frontend_0_n_115_12), .A1(
      frontend_0_n_115_2), .A2(frontend_0_n_120), .B1(inst_type[2]), .B2(
      frontend_0_n_190));
  INV_X1_LVT frontend_0_i_115_21 (.ZN(inst_src[8]), .A(frontend_0_n_115_12));
  INV_X1_LVT frontend_0_i_114_7 (.ZN(frontend_0_n_114_7), .A(
      frontend_0_inst_src_bin[3]));
  NAND2_X1_LVT frontend_0_i_114_9 (.ZN(frontend_0_n_114_9), .A1(
      frontend_0_inst_src_bin[2]), .A2(frontend_0_n_114_7));
  NOR2_X1_LVT frontend_0_i_114_19 (.ZN(frontend_0_n_189), .A1(frontend_0_n_114_5), 
      .A2(frontend_0_n_114_9));
  AOI22_X1_LVT frontend_0_i_115_18 (.ZN(frontend_0_n_115_11), .A1(
      frontend_0_n_115_2), .A2(frontend_0_n_119), .B1(inst_type[2]), .B2(
      frontend_0_n_189));
  INV_X1_LVT frontend_0_i_115_19 (.ZN(inst_src[7]), .A(frontend_0_n_115_11));
  NOR2_X1_LVT frontend_0_i_114_18 (.ZN(frontend_0_n_188), .A1(frontend_0_n_114_4), 
      .A2(frontend_0_n_114_9));
  AOI22_X1_LVT frontend_0_i_115_16 (.ZN(frontend_0_n_115_10), .A1(
      frontend_0_n_115_2), .A2(frontend_0_n_118), .B1(inst_type[2]), .B2(
      frontend_0_n_188));
  INV_X1_LVT frontend_0_i_115_17 (.ZN(inst_src[6]), .A(frontend_0_n_115_10));
  NOR2_X1_LVT frontend_0_i_114_17 (.ZN(frontend_0_n_187), .A1(frontend_0_n_114_3), 
      .A2(frontend_0_n_114_9));
  AOI22_X1_LVT frontend_0_i_115_14 (.ZN(frontend_0_n_115_9), .A1(
      frontend_0_n_115_2), .A2(frontend_0_n_117), .B1(inst_type[2]), .B2(
      frontend_0_n_187));
  INV_X1_LVT frontend_0_i_115_15 (.ZN(inst_src[5]), .A(frontend_0_n_115_9));
  NOR2_X1_LVT frontend_0_i_114_16 (.ZN(frontend_0_n_186), .A1(frontend_0_n_114_2), 
      .A2(frontend_0_n_114_9));
  AOI22_X1_LVT frontend_0_i_115_12 (.ZN(frontend_0_n_115_8), .A1(
      frontend_0_n_115_2), .A2(frontend_0_n_116), .B1(inst_type[2]), .B2(
      frontend_0_n_186));
  INV_X1_LVT frontend_0_i_115_13 (.ZN(inst_src[4]), .A(frontend_0_n_115_8));
  NAND2_X1_LVT frontend_0_i_114_8 (.ZN(frontend_0_n_114_8), .A1(
      frontend_0_n_114_6), .A2(frontend_0_n_114_7));
  NOR2_X1_LVT frontend_0_i_114_15 (.ZN(frontend_0_n_185), .A1(frontend_0_n_114_5), 
      .A2(frontend_0_n_114_8));
  AOI22_X1_LVT frontend_0_i_115_10 (.ZN(frontend_0_n_115_7), .A1(
      frontend_0_n_115_2), .A2(frontend_0_n_115), .B1(inst_type[2]), .B2(
      frontend_0_n_185));
  INV_X1_LVT frontend_0_i_115_11 (.ZN(inst_src[3]), .A(frontend_0_n_115_7));
  NOR2_X1_LVT frontend_0_i_114_14 (.ZN(frontend_0_n_184), .A1(frontend_0_n_114_4), 
      .A2(frontend_0_n_114_8));
  AOI22_X1_LVT frontend_0_i_115_8 (.ZN(frontend_0_n_115_6), .A1(
      frontend_0_n_115_2), .A2(frontend_0_n_114), .B1(inst_type[2]), .B2(
      frontend_0_n_184));
  INV_X1_LVT frontend_0_i_115_9 (.ZN(inst_src[2]), .A(frontend_0_n_115_6));
  INV_X1_LVT frontend_0_i_115_5 (.ZN(frontend_0_n_115_4), .A(inst_type[2]));
  NOR2_X1_LVT frontend_0_i_114_13 (.ZN(frontend_0_n_183), .A1(frontend_0_n_114_3), 
      .A2(frontend_0_n_114_8));
  AOI222_X1_LVT frontend_0_i_115_6 (.ZN(frontend_0_n_115_5), .A1(
      frontend_0_n_115_2), .A2(frontend_0_n_113), .B1(frontend_0_n_115_4), .B2(
      inst_so[6]), .C1(inst_type[2]), .C2(frontend_0_n_183));
  INV_X1_LVT frontend_0_i_115_7 (.ZN(inst_src[1]), .A(frontend_0_n_115_5));
  NOR2_X1_LVT frontend_0_i_114_12 (.ZN(frontend_0_n_182), .A1(frontend_0_n_114_2), 
      .A2(frontend_0_n_114_8));
  AOI222_X1_LVT frontend_0_i_115_3 (.ZN(frontend_0_n_115_3), .A1(
      frontend_0_n_115_2), .A2(frontend_0_n_112), .B1(frontend_0_n_115_0), .B2(
      inst_so[7]), .C1(frontend_0_n_182), .C2(inst_type[2]));
  INV_X1_LVT frontend_0_i_115_4 (.ZN(inst_src[0]), .A(frontend_0_n_115_3));
  NOR3_X1_LVT frontend_0_i_6_7 (.ZN(frontend_0_n_8), .A1(frontend_0_i_state[0]), 
      .A2(frontend_0_i_state[1]), .A3(frontend_0_i_state[2]));
  NOR2_X1_LVT frontend_0_i_118_0 (.ZN(frontend_0_n_118_0), .A1(irq[13]), .A2(
      nmi_pnd));
  INV_X1_LVT frontend_0_i_118_1 (.ZN(frontend_0_n_118_1), .A(frontend_0_n_118_0));
  NOR2_X1_LVT frontend_0_i_118_2 (.ZN(frontend_0_n_118_2), .A1(
      frontend_0_n_118_1), .A2(irq[12]));
  INV_X1_LVT frontend_0_i_118_3 (.ZN(frontend_0_n_118_3), .A(frontend_0_n_118_2));
  NOR2_X1_LVT frontend_0_i_118_4 (.ZN(frontend_0_n_118_4), .A1(
      frontend_0_n_118_3), .A2(irq[11]));
  INV_X1_LVT frontend_0_i_118_5 (.ZN(frontend_0_n_118_5), .A(frontend_0_n_118_4));
  OR2_X1_LVT frontend_0_i_116_0 (.ZN(frontend_0_n_198), .A1(irq[10]), .A2(
      wdt_irq));
  NOR2_X1_LVT frontend_0_i_118_6 (.ZN(frontend_0_n_118_6), .A1(
      frontend_0_n_118_5), .A2(frontend_0_n_198));
  INV_X1_LVT frontend_0_i_118_7 (.ZN(frontend_0_n_118_7), .A(irq[9]));
  NAND2_X1_LVT frontend_0_i_118_8 (.ZN(frontend_0_n_118_8), .A1(
      frontend_0_n_118_6), .A2(frontend_0_n_118_7));
  NOR2_X1_LVT frontend_0_i_118_9 (.ZN(frontend_0_n_118_9), .A1(
      frontend_0_n_118_8), .A2(irq[8]));
  INV_X1_LVT frontend_0_i_118_10 (.ZN(frontend_0_n_118_10), .A(
      frontend_0_n_118_9));
  NOR2_X1_LVT frontend_0_i_118_11 (.ZN(frontend_0_n_118_11), .A1(
      frontend_0_n_118_10), .A2(irq[7]));
  INV_X1_LVT frontend_0_i_118_12 (.ZN(frontend_0_n_118_12), .A(
      frontend_0_n_118_11));
  NOR2_X1_LVT frontend_0_i_118_13 (.ZN(frontend_0_n_118_13), .A1(
      frontend_0_n_118_12), .A2(irq[6]));
  INV_X1_LVT frontend_0_i_118_14 (.ZN(frontend_0_n_118_14), .A(irq[5]));
  NAND2_X1_LVT frontend_0_i_118_15 (.ZN(frontend_0_n_118_15), .A1(
      frontend_0_n_118_13), .A2(frontend_0_n_118_14));
  NOR2_X1_LVT frontend_0_i_118_16 (.ZN(frontend_0_n_118_16), .A1(
      frontend_0_n_118_15), .A2(irq[4]));
  INV_X1_LVT frontend_0_i_118_17 (.ZN(frontend_0_n_118_17), .A(irq[3]));
  NAND2_X1_LVT frontend_0_i_118_18 (.ZN(frontend_0_n_118_18), .A1(
      frontend_0_n_118_16), .A2(frontend_0_n_118_17));
  NOR2_X1_LVT frontend_0_i_118_19 (.ZN(frontend_0_n_118_19), .A1(
      frontend_0_n_118_18), .A2(irq[2]));
  NAND2_X1_LVT frontend_0_i_118_20 (.ZN(frontend_0_n_118_20), .A1(
      frontend_0_n_118_19), .A2(irq[1]));
  INV_X1_LVT frontend_0_i_118_21 (.ZN(frontend_0_n_118_21), .A(
      frontend_0_n_118_20));
  NAND2_X1_LVT frontend_0_i_118_22 (.ZN(frontend_0_n_118_22), .A1(
      frontend_0_n_118_9), .A2(irq[7]));
  NAND2_X1_LVT frontend_0_i_118_23 (.ZN(frontend_0_n_118_23), .A1(
      frontend_0_n_118_6), .A2(irq[9]));
  NAND2_X1_LVT frontend_0_i_118_24 (.ZN(frontend_0_n_118_24), .A1(
      frontend_0_n_118_2), .A2(irq[11]));
  INV_X1_LVT frontend_0_i_118_25 (.ZN(frontend_0_n_118_25), .A(nmi_pnd));
  NAND2_X1_LVT frontend_0_i_118_26 (.ZN(frontend_0_n_118_26), .A1(
      frontend_0_n_118_25), .A2(irq[13]));
  NAND4_X1_LVT frontend_0_i_118_27 (.ZN(frontend_0_n_118_27), .A1(
      frontend_0_n_118_22), .A2(frontend_0_n_118_23), .A3(frontend_0_n_118_24), 
      .A4(frontend_0_n_118_26));
  AND2_X1_LVT frontend_0_i_118_28 (.ZN(frontend_0_n_118_28), .A1(
      frontend_0_n_118_16), .A2(irq[3]));
  NAND2_X1_LVT frontend_0_i_118_29 (.ZN(frontend_0_n_118_29), .A1(
      frontend_0_n_118_13), .A2(irq[5]));
  INV_X1_LVT frontend_0_i_118_30 (.ZN(frontend_0_n_118_30), .A(
      frontend_0_n_118_29));
  NOR4_X1_LVT frontend_0_i_118_31 (.ZN(frontend_0_n_118_31), .A1(
      frontend_0_n_118_21), .A2(frontend_0_n_118_27), .A3(frontend_0_n_118_28), 
      .A4(frontend_0_n_118_30));
  INV_X1_LVT frontend_0_i_118_32 (.ZN(frontend_0_n_118_32), .A(
      frontend_0_n_118_19));
  NOR2_X1_LVT frontend_0_i_118_33 (.ZN(frontend_0_n_118_33), .A1(
      frontend_0_n_118_32), .A2(irq[1]));
  INV_X1_LVT frontend_0_i_118_34 (.ZN(frontend_0_n_118_34), .A(irq[0]));
  NAND2_X1_LVT frontend_0_i_118_35 (.ZN(frontend_0_n_118_35), .A1(
      frontend_0_n_118_33), .A2(frontend_0_n_118_34));
  NAND2_X1_LVT frontend_0_i_118_36 (.ZN(frontend_0_n_200), .A1(
      frontend_0_n_118_31), .A2(frontend_0_n_118_35));
  CLKGATETST_X1_LVT frontend_0_clk_gate_irq_num_reg (.GCK(frontend_0_n_199), .CK(
      cpu_mclk), .E(frontend_0_irq_detect), .SE(1'b0));
  DFFS_X1_LVT \frontend_0_irq_num_reg[0] (.Q(frontend_0_irq_num[0]), .QN(), .CK(
      frontend_0_n_199), .D(frontend_0_n_200), .SN(frontend_0_n_91));
  INV_X1_LVT frontend_0_i_120_0 (.ZN(frontend_0_n_120_0), .A(
      frontend_0_irq_num[0]));
  INV_X1_LVT frontend_0_i_118_37 (.ZN(frontend_0_n_118_36), .A(irq[2]));
  NOR2_X1_LVT frontend_0_i_118_38 (.ZN(frontend_0_n_118_37), .A1(
      frontend_0_n_118_18), .A2(frontend_0_n_118_36));
  NAND2_X1_LVT frontend_0_i_118_39 (.ZN(frontend_0_n_118_38), .A1(
      frontend_0_n_118_4), .A2(frontend_0_n_198));
  NAND4_X1_LVT frontend_0_i_118_40 (.ZN(frontend_0_n_118_39), .A1(
      frontend_0_n_118_22), .A2(frontend_0_n_118_38), .A3(frontend_0_n_118_24), 
      .A4(frontend_0_n_118_25));
  NAND2_X1_LVT frontend_0_i_118_41 (.ZN(frontend_0_n_118_40), .A1(
      frontend_0_n_118_11), .A2(irq[6]));
  INV_X1_LVT frontend_0_i_118_42 (.ZN(frontend_0_n_118_41), .A(
      frontend_0_n_118_40));
  NOR4_X1_LVT frontend_0_i_118_43 (.ZN(frontend_0_n_118_42), .A1(
      frontend_0_n_118_37), .A2(frontend_0_n_118_39), .A3(frontend_0_n_118_28), 
      .A4(frontend_0_n_118_41));
  NAND2_X1_LVT frontend_0_i_118_44 (.ZN(frontend_0_n_201), .A1(
      frontend_0_n_118_42), .A2(frontend_0_n_118_35));
  DFFS_X1_LVT \frontend_0_irq_num_reg[1] (.Q(frontend_0_irq_num[1]), .QN(), .CK(
      frontend_0_n_199), .D(frontend_0_n_201), .SN(frontend_0_n_91));
  NOR2_X1_LVT frontend_0_i_120_3 (.ZN(frontend_0_n_120_3), .A1(
      frontend_0_n_120_0), .A2(frontend_0_irq_num[1]));
  NAND2_X1_LVT frontend_0_i_118_45 (.ZN(frontend_0_n_118_43), .A1(
      frontend_0_n_118_0), .A2(irq[12]));
  NAND4_X1_LVT frontend_0_i_118_46 (.ZN(frontend_0_n_118_44), .A1(
      frontend_0_n_118_22), .A2(frontend_0_n_118_43), .A3(frontend_0_n_118_26), 
      .A4(frontend_0_n_118_25));
  INV_X1_LVT frontend_0_i_118_47 (.ZN(frontend_0_n_118_45), .A(irq[4]));
  NOR2_X1_LVT frontend_0_i_118_48 (.ZN(frontend_0_n_118_46), .A1(
      frontend_0_n_118_15), .A2(frontend_0_n_118_45));
  NOR4_X1_LVT frontend_0_i_118_49 (.ZN(frontend_0_n_118_47), .A1(
      frontend_0_n_118_44), .A2(frontend_0_n_118_46), .A3(frontend_0_n_118_30), 
      .A4(frontend_0_n_118_41));
  NAND2_X1_LVT frontend_0_i_118_50 (.ZN(frontend_0_n_202), .A1(
      frontend_0_n_118_47), .A2(frontend_0_n_118_35));
  DFFS_X1_LVT \frontend_0_irq_num_reg[2] (.Q(frontend_0_irq_num[2]), .QN(), .CK(
      frontend_0_n_199), .D(frontend_0_n_202), .SN(frontend_0_n_91));
  NAND2_X1_LVT frontend_0_i_120_12 (.ZN(frontend_0_n_120_12), .A1(
      frontend_0_n_120_3), .A2(frontend_0_irq_num[2]));
  NAND4_X1_LVT frontend_0_i_118_51 (.ZN(frontend_0_n_118_48), .A1(
      frontend_0_n_118_24), .A2(frontend_0_n_118_43), .A3(frontend_0_n_118_26), 
      .A4(frontend_0_n_118_25));
  INV_X1_LVT frontend_0_i_118_52 (.ZN(frontend_0_n_118_49), .A(irq[8]));
  NOR2_X1_LVT frontend_0_i_118_53 (.ZN(frontend_0_n_118_50), .A1(
      frontend_0_n_118_8), .A2(frontend_0_n_118_49));
  INV_X1_LVT frontend_0_i_118_54 (.ZN(frontend_0_n_118_51), .A(
      frontend_0_n_118_23));
  INV_X1_LVT frontend_0_i_118_55 (.ZN(frontend_0_n_118_52), .A(
      frontend_0_n_118_38));
  NOR4_X1_LVT frontend_0_i_118_56 (.ZN(frontend_0_n_118_53), .A1(
      frontend_0_n_118_48), .A2(frontend_0_n_118_50), .A3(frontend_0_n_118_51), 
      .A4(frontend_0_n_118_52));
  NAND2_X1_LVT frontend_0_i_118_57 (.ZN(frontend_0_n_203), .A1(
      frontend_0_n_118_53), .A2(frontend_0_n_118_35));
  DFFS_X1_LVT \frontend_0_irq_num_reg[3] (.Q(frontend_0_irq_num[3]), .QN(), .CK(
      frontend_0_n_199), .D(frontend_0_n_203), .SN(frontend_0_n_91));
  INV_X1_LVT frontend_0_i_120_15 (.ZN(frontend_0_n_120_15), .A(
      frontend_0_irq_num[3]));
  NAND4_X1_LVT frontend_0_i_118_58 (.ZN(frontend_0_n_118_54), .A1(
      frontend_0_n_118_53), .A2(frontend_0_n_118_29), .A3(frontend_0_n_118_40), 
      .A4(frontend_0_n_118_22));
  NOR4_X1_LVT frontend_0_i_118_59 (.ZN(frontend_0_n_118_55), .A1(
      frontend_0_n_118_54), .A2(frontend_0_n_118_37), .A3(frontend_0_n_118_28), 
      .A4(frontend_0_n_118_46));
  NAND2_X1_LVT frontend_0_i_118_60 (.ZN(frontend_0_n_118_56), .A1(
      frontend_0_n_118_33), .A2(irq[0]));
  NAND4_X1_LVT frontend_0_i_118_61 (.ZN(frontend_0_n_204), .A1(
      frontend_0_n_118_55), .A2(frontend_0_n_118_56), .A3(frontend_0_n_118_35), 
      .A4(frontend_0_n_118_20));
  DFFS_X1_LVT \frontend_0_irq_num_reg[4] (.Q(frontend_0_irq_num[4]), .QN(), .CK(
      frontend_0_n_199), .D(frontend_0_n_204), .SN(frontend_0_n_91));
  INV_X1_LVT frontend_0_i_120_16 (.ZN(frontend_0_n_120_16), .A(
      frontend_0_irq_num[4]));
  NOR2_X1_LVT frontend_0_i_120_18 (.ZN(frontend_0_n_120_18), .A1(
      frontend_0_n_120_15), .A2(frontend_0_n_120_16));
  DFFS_X1_LVT \frontend_0_irq_num_reg[5] (.Q(frontend_0_irq_num[5]), .QN(), .CK(
      frontend_0_n_199), .D(frontend_0_n_204), .SN(frontend_0_n_91));
  NAND2_X1_LVT frontend_0_i_120_20 (.ZN(frontend_0_n_120_20), .A1(
      frontend_0_n_120_18), .A2(frontend_0_irq_num[5]));
  NOR2_X1_LVT frontend_0_i_120_34 (.ZN(frontend_0_n_218), .A1(
      frontend_0_n_120_12), .A2(frontend_0_n_120_20));
  AND2_X1_LVT frontend_0_i_121_13 (.ZN(irq_acc[13]), .A1(frontend_0_n_8), .A2(
      frontend_0_n_218));
  NOR2_X1_LVT frontend_0_i_120_2 (.ZN(frontend_0_n_120_2), .A1(
      frontend_0_irq_num[0]), .A2(frontend_0_irq_num[1]));
  NAND2_X1_LVT frontend_0_i_120_11 (.ZN(frontend_0_n_120_11), .A1(
      frontend_0_n_120_2), .A2(frontend_0_irq_num[2]));
  NOR2_X1_LVT frontend_0_i_120_33 (.ZN(frontend_0_n_217), .A1(
      frontend_0_n_120_11), .A2(frontend_0_n_120_20));
  AND2_X1_LVT frontend_0_i_121_12 (.ZN(irq_acc[12]), .A1(frontend_0_n_8), .A2(
      frontend_0_n_217));
  INV_X1_LVT frontend_0_i_120_1 (.ZN(frontend_0_n_120_1), .A(
      frontend_0_irq_num[1]));
  NOR2_X1_LVT frontend_0_i_120_5 (.ZN(frontend_0_n_120_5), .A1(
      frontend_0_n_120_0), .A2(frontend_0_n_120_1));
  INV_X1_LVT frontend_0_i_120_6 (.ZN(frontend_0_n_120_6), .A(
      frontend_0_irq_num[2]));
  NAND2_X1_LVT frontend_0_i_120_10 (.ZN(frontend_0_n_120_10), .A1(
      frontend_0_n_120_5), .A2(frontend_0_n_120_6));
  NOR2_X1_LVT frontend_0_i_120_32 (.ZN(frontend_0_n_216), .A1(
      frontend_0_n_120_10), .A2(frontend_0_n_120_20));
  AND2_X1_LVT frontend_0_i_121_11 (.ZN(irq_acc[11]), .A1(frontend_0_n_8), .A2(
      frontend_0_n_216));
  NOR2_X1_LVT frontend_0_i_120_4 (.ZN(frontend_0_n_120_4), .A1(
      frontend_0_irq_num[0]), .A2(frontend_0_n_120_1));
  NAND2_X1_LVT frontend_0_i_120_9 (.ZN(frontend_0_n_120_9), .A1(
      frontend_0_n_120_4), .A2(frontend_0_n_120_6));
  NOR2_X1_LVT frontend_0_i_120_31 (.ZN(frontend_0_n_215), .A1(frontend_0_n_120_9), 
      .A2(frontend_0_n_120_20));
  AND2_X1_LVT frontend_0_i_121_10 (.ZN(irq_acc[10]), .A1(frontend_0_n_8), .A2(
      frontend_0_n_215));
  NAND2_X1_LVT frontend_0_i_120_8 (.ZN(frontend_0_n_120_8), .A1(
      frontend_0_n_120_3), .A2(frontend_0_n_120_6));
  NOR2_X1_LVT frontend_0_i_120_30 (.ZN(frontend_0_n_214), .A1(frontend_0_n_120_8), 
      .A2(frontend_0_n_120_20));
  AND2_X1_LVT frontend_0_i_121_9 (.ZN(irq_acc[9]), .A1(frontend_0_n_8), .A2(
      frontend_0_n_214));
  NAND2_X1_LVT frontend_0_i_120_7 (.ZN(frontend_0_n_120_7), .A1(
      frontend_0_n_120_2), .A2(frontend_0_n_120_6));
  NOR2_X1_LVT frontend_0_i_120_29 (.ZN(frontend_0_n_213), .A1(frontend_0_n_120_7), 
      .A2(frontend_0_n_120_20));
  AND2_X1_LVT frontend_0_i_121_8 (.ZN(irq_acc[8]), .A1(frontend_0_n_8), .A2(
      frontend_0_n_213));
  NAND2_X1_LVT frontend_0_i_120_14 (.ZN(frontend_0_n_120_14), .A1(
      frontend_0_n_120_5), .A2(frontend_0_irq_num[2]));
  NOR2_X1_LVT frontend_0_i_120_17 (.ZN(frontend_0_n_120_17), .A1(
      frontend_0_irq_num[3]), .A2(frontend_0_n_120_16));
  NAND2_X1_LVT frontend_0_i_120_19 (.ZN(frontend_0_n_120_19), .A1(
      frontend_0_n_120_17), .A2(frontend_0_irq_num[5]));
  NOR2_X1_LVT frontend_0_i_120_28 (.ZN(frontend_0_n_212), .A1(
      frontend_0_n_120_14), .A2(frontend_0_n_120_19));
  AND2_X1_LVT frontend_0_i_121_7 (.ZN(irq_acc[7]), .A1(frontend_0_n_8), .A2(
      frontend_0_n_212));
  NAND2_X1_LVT frontend_0_i_120_13 (.ZN(frontend_0_n_120_13), .A1(
      frontend_0_n_120_4), .A2(frontend_0_irq_num[2]));
  NOR2_X1_LVT frontend_0_i_120_27 (.ZN(frontend_0_n_211), .A1(
      frontend_0_n_120_13), .A2(frontend_0_n_120_19));
  AND2_X1_LVT frontend_0_i_121_6 (.ZN(irq_acc[6]), .A1(frontend_0_n_8), .A2(
      frontend_0_n_211));
  NOR2_X1_LVT frontend_0_i_120_26 (.ZN(frontend_0_n_210), .A1(
      frontend_0_n_120_12), .A2(frontend_0_n_120_19));
  AND2_X1_LVT frontend_0_i_121_5 (.ZN(irq_acc[5]), .A1(frontend_0_n_8), .A2(
      frontend_0_n_210));
  NOR2_X1_LVT frontend_0_i_120_25 (.ZN(frontend_0_n_209), .A1(
      frontend_0_n_120_11), .A2(frontend_0_n_120_19));
  AND2_X1_LVT frontend_0_i_121_4 (.ZN(irq_acc[4]), .A1(frontend_0_n_8), .A2(
      frontend_0_n_209));
  NOR2_X1_LVT frontend_0_i_120_24 (.ZN(frontend_0_n_208), .A1(
      frontend_0_n_120_10), .A2(frontend_0_n_120_19));
  AND2_X1_LVT frontend_0_i_121_3 (.ZN(irq_acc[3]), .A1(frontend_0_n_8), .A2(
      frontend_0_n_208));
  NOR2_X1_LVT frontend_0_i_120_23 (.ZN(frontend_0_n_207), .A1(frontend_0_n_120_9), 
      .A2(frontend_0_n_120_19));
  AND2_X1_LVT frontend_0_i_121_2 (.ZN(irq_acc[2]), .A1(frontend_0_n_8), .A2(
      frontend_0_n_207));
  NOR2_X1_LVT frontend_0_i_120_22 (.ZN(frontend_0_n_206), .A1(frontend_0_n_120_8), 
      .A2(frontend_0_n_120_19));
  AND2_X1_LVT frontend_0_i_121_1 (.ZN(irq_acc[1]), .A1(frontend_0_n_8), .A2(
      frontend_0_n_206));
  NOR2_X1_LVT frontend_0_i_120_21 (.ZN(frontend_0_n_205), .A1(frontend_0_n_120_7), 
      .A2(frontend_0_n_120_19));
  AND2_X1_LVT frontend_0_i_121_0 (.ZN(irq_acc[0]), .A1(frontend_0_n_8), .A2(
      frontend_0_n_205));
  INV_X1_LVT frontend_0_i_127_0 (.ZN(frontend_0_n_127_0), .A(pc_sw_wr));
  NOR3_X1_LVT frontend_0_i_125_2 (.ZN(frontend_0_n_221), .A1(
      frontend_0_i_state[0]), .A2(frontend_0_i_state[1]), .A3(
      frontend_0_i_state[2]));
  INV_X1_LVT frontend_0_i_125_0 (.ZN(frontend_0_n_125_0), .A(
      frontend_0_i_state[0]));
  NOR3_X1_LVT frontend_0_i_125_1 (.ZN(frontend_0_n_220), .A1(frontend_0_n_125_0), 
      .A2(frontend_0_i_state[1]), .A3(frontend_0_i_state[2]));
  NOR2_X1_LVT frontend_0_i_125_3 (.ZN(frontend_0_n_222), .A1(frontend_0_n_220), 
      .A2(frontend_0_n_221));
  DFFR_X1_LVT \frontend_0_pc_reg[15] (.Q(pc[15]), .QN(), .CK(cpu_mclk), .D(
      pc_nxt[15]), .RN(frontend_0_n_91));
  AOI221_X1_LVT frontend_0_i_126_28 (.ZN(frontend_0_n_126_14), .A(
      frontend_0_n_221), .B1(frontend_0_n_220), .B2(fe_mdb_in[14]), .C1(
      frontend_0_n_222), .C2(frontend_0_pc_incr[14]));
  INV_X1_LVT frontend_0_i_126_29 (.ZN(frontend_0_n_237), .A(frontend_0_n_126_14));
  AOI22_X1_LVT frontend_0_i_127_29 (.ZN(frontend_0_n_127_15), .A1(
      frontend_0_n_127_0), .A2(frontend_0_n_237), .B1(pc_sw_wr), .B2(pc_sw[14]));
  INV_X1_LVT frontend_0_i_127_30 (.ZN(pc_nxt[14]), .A(frontend_0_n_127_15));
  DFFR_X1_LVT \frontend_0_pc_reg[14] (.Q(pc[14]), .QN(), .CK(cpu_mclk), .D(
      pc_nxt[14]), .RN(frontend_0_n_91));
  AOI221_X1_LVT frontend_0_i_126_26 (.ZN(frontend_0_n_126_13), .A(
      frontend_0_n_221), .B1(frontend_0_n_220), .B2(fe_mdb_in[13]), .C1(
      frontend_0_n_222), .C2(frontend_0_pc_incr[13]));
  INV_X1_LVT frontend_0_i_126_27 (.ZN(frontend_0_n_236), .A(frontend_0_n_126_13));
  AOI22_X1_LVT frontend_0_i_127_27 (.ZN(frontend_0_n_127_14), .A1(
      frontend_0_n_127_0), .A2(frontend_0_n_236), .B1(pc_sw_wr), .B2(pc_sw[13]));
  INV_X1_LVT frontend_0_i_127_28 (.ZN(pc_nxt[13]), .A(frontend_0_n_127_14));
  DFFR_X1_LVT \frontend_0_pc_reg[13] (.Q(pc[13]), .QN(), .CK(cpu_mclk), .D(
      pc_nxt[13]), .RN(frontend_0_n_91));
  AOI221_X1_LVT frontend_0_i_126_24 (.ZN(frontend_0_n_126_12), .A(
      frontend_0_n_221), .B1(frontend_0_n_220), .B2(fe_mdb_in[12]), .C1(
      frontend_0_n_222), .C2(frontend_0_pc_incr[12]));
  INV_X1_LVT frontend_0_i_126_25 (.ZN(frontend_0_n_235), .A(frontend_0_n_126_12));
  AOI22_X1_LVT frontend_0_i_127_25 (.ZN(frontend_0_n_127_13), .A1(
      frontend_0_n_127_0), .A2(frontend_0_n_235), .B1(pc_sw_wr), .B2(pc_sw[12]));
  INV_X1_LVT frontend_0_i_127_26 (.ZN(pc_nxt[12]), .A(frontend_0_n_127_13));
  DFFR_X1_LVT \frontend_0_pc_reg[12] (.Q(pc[12]), .QN(), .CK(cpu_mclk), .D(
      pc_nxt[12]), .RN(frontend_0_n_91));
  AOI221_X1_LVT frontend_0_i_126_22 (.ZN(frontend_0_n_126_11), .A(
      frontend_0_n_221), .B1(frontend_0_n_220), .B2(fe_mdb_in[11]), .C1(
      frontend_0_n_222), .C2(frontend_0_pc_incr[11]));
  INV_X1_LVT frontend_0_i_126_23 (.ZN(frontend_0_n_234), .A(frontend_0_n_126_11));
  AOI22_X1_LVT frontend_0_i_127_23 (.ZN(frontend_0_n_127_12), .A1(
      frontend_0_n_127_0), .A2(frontend_0_n_234), .B1(pc_sw_wr), .B2(pc_sw[11]));
  INV_X1_LVT frontend_0_i_127_24 (.ZN(pc_nxt[11]), .A(frontend_0_n_127_12));
  DFFR_X1_LVT \frontend_0_pc_reg[11] (.Q(pc[11]), .QN(), .CK(cpu_mclk), .D(
      pc_nxt[11]), .RN(frontend_0_n_91));
  AOI221_X1_LVT frontend_0_i_126_20 (.ZN(frontend_0_n_126_10), .A(
      frontend_0_n_221), .B1(frontend_0_n_220), .B2(fe_mdb_in[10]), .C1(
      frontend_0_n_222), .C2(frontend_0_pc_incr[10]));
  INV_X1_LVT frontend_0_i_126_21 (.ZN(frontend_0_n_233), .A(frontend_0_n_126_10));
  AOI22_X1_LVT frontend_0_i_127_21 (.ZN(frontend_0_n_127_11), .A1(
      frontend_0_n_127_0), .A2(frontend_0_n_233), .B1(pc_sw_wr), .B2(pc_sw[10]));
  INV_X1_LVT frontend_0_i_127_22 (.ZN(pc_nxt[10]), .A(frontend_0_n_127_11));
  DFFR_X1_LVT \frontend_0_pc_reg[10] (.Q(pc[10]), .QN(), .CK(cpu_mclk), .D(
      pc_nxt[10]), .RN(frontend_0_n_91));
  AOI221_X1_LVT frontend_0_i_126_18 (.ZN(frontend_0_n_126_9), .A(
      frontend_0_n_221), .B1(frontend_0_n_220), .B2(fe_mdb_in[9]), .C1(
      frontend_0_n_222), .C2(frontend_0_pc_incr[9]));
  INV_X1_LVT frontend_0_i_126_19 (.ZN(frontend_0_n_232), .A(frontend_0_n_126_9));
  AOI22_X1_LVT frontend_0_i_127_19 (.ZN(frontend_0_n_127_10), .A1(
      frontend_0_n_127_0), .A2(frontend_0_n_232), .B1(pc_sw_wr), .B2(pc_sw[9]));
  INV_X1_LVT frontend_0_i_127_20 (.ZN(pc_nxt[9]), .A(frontend_0_n_127_10));
  DFFR_X1_LVT \frontend_0_pc_reg[9] (.Q(pc[9]), .QN(), .CK(cpu_mclk), .D(
      pc_nxt[9]), .RN(frontend_0_n_91));
  AOI221_X1_LVT frontend_0_i_126_16 (.ZN(frontend_0_n_126_8), .A(
      frontend_0_n_221), .B1(frontend_0_n_220), .B2(fe_mdb_in[8]), .C1(
      frontend_0_n_222), .C2(frontend_0_pc_incr[8]));
  INV_X1_LVT frontend_0_i_126_17 (.ZN(frontend_0_n_231), .A(frontend_0_n_126_8));
  AOI22_X1_LVT frontend_0_i_127_17 (.ZN(frontend_0_n_127_9), .A1(
      frontend_0_n_127_0), .A2(frontend_0_n_231), .B1(pc_sw_wr), .B2(pc_sw[8]));
  INV_X1_LVT frontend_0_i_127_18 (.ZN(pc_nxt[8]), .A(frontend_0_n_127_9));
  DFFR_X1_LVT \frontend_0_pc_reg[8] (.Q(pc[8]), .QN(), .CK(cpu_mclk), .D(
      pc_nxt[8]), .RN(frontend_0_n_91));
  AOI221_X1_LVT frontend_0_i_126_14 (.ZN(frontend_0_n_126_7), .A(
      frontend_0_n_221), .B1(frontend_0_n_220), .B2(fe_mdb_in[7]), .C1(
      frontend_0_n_222), .C2(frontend_0_pc_incr[7]));
  INV_X1_LVT frontend_0_i_126_15 (.ZN(frontend_0_n_230), .A(frontend_0_n_126_7));
  AOI22_X1_LVT frontend_0_i_127_15 (.ZN(frontend_0_n_127_8), .A1(
      frontend_0_n_127_0), .A2(frontend_0_n_230), .B1(pc_sw_wr), .B2(pc_sw[7]));
  INV_X1_LVT frontend_0_i_127_16 (.ZN(pc_nxt[7]), .A(frontend_0_n_127_8));
  DFFR_X1_LVT \frontend_0_pc_reg[7] (.Q(pc[7]), .QN(), .CK(cpu_mclk), .D(
      pc_nxt[7]), .RN(frontend_0_n_91));
  AOI222_X1_LVT frontend_0_i_126_12 (.ZN(frontend_0_n_126_6), .A1(
      frontend_0_n_221), .A2(frontend_0_irq_num[5]), .B1(frontend_0_n_220), .B2(
      fe_mdb_in[6]), .C1(frontend_0_n_222), .C2(frontend_0_pc_incr[6]));
  INV_X1_LVT frontend_0_i_126_13 (.ZN(frontend_0_n_229), .A(frontend_0_n_126_6));
  AOI22_X1_LVT frontend_0_i_127_13 (.ZN(frontend_0_n_127_7), .A1(
      frontend_0_n_127_0), .A2(frontend_0_n_229), .B1(pc_sw_wr), .B2(pc_sw[6]));
  INV_X1_LVT frontend_0_i_127_14 (.ZN(pc_nxt[6]), .A(frontend_0_n_127_7));
  DFFR_X1_LVT \frontend_0_pc_reg[6] (.Q(pc[6]), .QN(), .CK(cpu_mclk), .D(
      pc_nxt[6]), .RN(frontend_0_n_91));
  AOI222_X1_LVT frontend_0_i_126_10 (.ZN(frontend_0_n_126_5), .A1(
      frontend_0_n_221), .A2(frontend_0_irq_num[4]), .B1(frontend_0_n_220), .B2(
      fe_mdb_in[5]), .C1(frontend_0_n_222), .C2(frontend_0_pc_incr[5]));
  INV_X1_LVT frontend_0_i_126_11 (.ZN(frontend_0_n_228), .A(frontend_0_n_126_5));
  AOI22_X1_LVT frontend_0_i_127_11 (.ZN(frontend_0_n_127_6), .A1(
      frontend_0_n_127_0), .A2(frontend_0_n_228), .B1(pc_sw_wr), .B2(pc_sw[5]));
  INV_X1_LVT frontend_0_i_127_12 (.ZN(pc_nxt[5]), .A(frontend_0_n_127_6));
  DFFR_X1_LVT \frontend_0_pc_reg[5] (.Q(pc[5]), .QN(), .CK(cpu_mclk), .D(
      pc_nxt[5]), .RN(frontend_0_n_91));
  AOI222_X1_LVT frontend_0_i_126_8 (.ZN(frontend_0_n_126_4), .A1(
      frontend_0_n_221), .A2(frontend_0_irq_num[3]), .B1(frontend_0_n_220), .B2(
      fe_mdb_in[4]), .C1(frontend_0_n_222), .C2(frontend_0_pc_incr[4]));
  INV_X1_LVT frontend_0_i_126_9 (.ZN(frontend_0_n_227), .A(frontend_0_n_126_4));
  AOI22_X1_LVT frontend_0_i_127_9 (.ZN(frontend_0_n_127_5), .A1(
      frontend_0_n_127_0), .A2(frontend_0_n_227), .B1(pc_sw_wr), .B2(pc_sw[4]));
  INV_X1_LVT frontend_0_i_127_10 (.ZN(pc_nxt[4]), .A(frontend_0_n_127_5));
  DFFR_X1_LVT \frontend_0_pc_reg[4] (.Q(pc[4]), .QN(), .CK(cpu_mclk), .D(
      pc_nxt[4]), .RN(frontend_0_n_91));
  AOI222_X1_LVT frontend_0_i_126_6 (.ZN(frontend_0_n_126_3), .A1(
      frontend_0_n_221), .A2(frontend_0_irq_num[2]), .B1(frontend_0_n_220), .B2(
      fe_mdb_in[3]), .C1(frontend_0_n_222), .C2(frontend_0_pc_incr[3]));
  INV_X1_LVT frontend_0_i_126_7 (.ZN(frontend_0_n_226), .A(frontend_0_n_126_3));
  AOI22_X1_LVT frontend_0_i_127_7 (.ZN(frontend_0_n_127_4), .A1(
      frontend_0_n_127_0), .A2(frontend_0_n_226), .B1(pc_sw_wr), .B2(pc_sw[3]));
  INV_X1_LVT frontend_0_i_127_8 (.ZN(pc_nxt[3]), .A(frontend_0_n_127_4));
  DFFR_X1_LVT \frontend_0_pc_reg[3] (.Q(pc[3]), .QN(), .CK(cpu_mclk), .D(
      pc_nxt[3]), .RN(frontend_0_n_91));
  AOI222_X1_LVT frontend_0_i_126_4 (.ZN(frontend_0_n_126_2), .A1(
      frontend_0_n_221), .A2(frontend_0_irq_num[1]), .B1(frontend_0_n_220), .B2(
      fe_mdb_in[2]), .C1(frontend_0_n_222), .C2(frontend_0_pc_incr[2]));
  INV_X1_LVT frontend_0_i_126_5 (.ZN(frontend_0_n_225), .A(frontend_0_n_126_2));
  AOI22_X1_LVT frontend_0_i_127_5 (.ZN(frontend_0_n_127_3), .A1(
      frontend_0_n_127_0), .A2(frontend_0_n_225), .B1(pc_sw_wr), .B2(pc_sw[2]));
  INV_X1_LVT frontend_0_i_127_6 (.ZN(pc_nxt[2]), .A(frontend_0_n_127_3));
  DFFR_X1_LVT \frontend_0_pc_reg[2] (.Q(pc[2]), .QN(), .CK(cpu_mclk), .D(
      pc_nxt[2]), .RN(frontend_0_n_91));
  INV_X1_LVT frontend_0_i_122_0 (.ZN(frontend_0_n_122_0), .A(
      frontend_0_e_state_nxt_reg[1]));
  AND4_X1_LVT frontend_0_i_122_1 (.ZN(frontend_0_n_122_1), .A1(
      frontend_0_n_122_0), .A2(frontend_0_e_state_nxt_reg[0]), .A3(
      frontend_0_e_state_nxt_reg[2]), .A4(frontend_0_e_state_nxt_reg[3]));
  INV_X1_LVT frontend_0_i_122_2 (.ZN(frontend_0_n_122_2), .A(frontend_0_n_73));
  AOI21_X1_LVT frontend_0_i_122_3 (.ZN(frontend_0_fetch), .A(frontend_0_n_122_1), 
      .B1(frontend_0_n_122_2), .B2(frontend_0_n_4));
  AOI222_X1_LVT frontend_0_i_126_2 (.ZN(frontend_0_n_126_1), .A1(
      frontend_0_n_221), .A2(frontend_0_irq_num[0]), .B1(frontend_0_n_220), .B2(
      fe_mdb_in[1]), .C1(frontend_0_n_222), .C2(frontend_0_pc_incr[1]));
  INV_X1_LVT frontend_0_i_126_3 (.ZN(frontend_0_n_224), .A(frontend_0_n_126_1));
  AOI22_X1_LVT frontend_0_i_127_3 (.ZN(frontend_0_n_127_2), .A1(
      frontend_0_n_127_0), .A2(frontend_0_n_224), .B1(pc_sw_wr), .B2(pc_sw[1]));
  INV_X1_LVT frontend_0_i_127_4 (.ZN(pc_nxt[1]), .A(frontend_0_n_127_2));
  DFFR_X1_LVT \frontend_0_pc_reg[1] (.Q(pc[1]), .QN(), .CK(cpu_mclk), .D(
      pc_nxt[1]), .RN(frontend_0_n_91));
  HA_X1_LVT frontend_0_i_124_0 (.CO(frontend_0_n_124_0), .S(
      frontend_0_pc_incr[1]), .A(frontend_0_fetch), .B(pc[1]));
  HA_X1_LVT frontend_0_i_124_1 (.CO(frontend_0_n_124_1), .S(
      frontend_0_pc_incr[2]), .A(pc[2]), .B(frontend_0_n_124_0));
  HA_X1_LVT frontend_0_i_124_2 (.CO(frontend_0_n_124_2), .S(
      frontend_0_pc_incr[3]), .A(pc[3]), .B(frontend_0_n_124_1));
  HA_X1_LVT frontend_0_i_124_3 (.CO(frontend_0_n_124_3), .S(
      frontend_0_pc_incr[4]), .A(pc[4]), .B(frontend_0_n_124_2));
  HA_X1_LVT frontend_0_i_124_4 (.CO(frontend_0_n_124_4), .S(
      frontend_0_pc_incr[5]), .A(pc[5]), .B(frontend_0_n_124_3));
  HA_X1_LVT frontend_0_i_124_5 (.CO(frontend_0_n_124_5), .S(
      frontend_0_pc_incr[6]), .A(pc[6]), .B(frontend_0_n_124_4));
  HA_X1_LVT frontend_0_i_124_6 (.CO(frontend_0_n_124_6), .S(
      frontend_0_pc_incr[7]), .A(pc[7]), .B(frontend_0_n_124_5));
  HA_X1_LVT frontend_0_i_124_7 (.CO(frontend_0_n_124_7), .S(
      frontend_0_pc_incr[8]), .A(pc[8]), .B(frontend_0_n_124_6));
  HA_X1_LVT frontend_0_i_124_8 (.CO(frontend_0_n_124_8), .S(
      frontend_0_pc_incr[9]), .A(pc[9]), .B(frontend_0_n_124_7));
  HA_X1_LVT frontend_0_i_124_9 (.CO(frontend_0_n_124_9), .S(
      frontend_0_pc_incr[10]), .A(pc[10]), .B(frontend_0_n_124_8));
  HA_X1_LVT frontend_0_i_124_10 (.CO(frontend_0_n_124_10), .S(
      frontend_0_pc_incr[11]), .A(pc[11]), .B(frontend_0_n_124_9));
  HA_X1_LVT frontend_0_i_124_11 (.CO(frontend_0_n_124_11), .S(
      frontend_0_pc_incr[12]), .A(pc[12]), .B(frontend_0_n_124_10));
  HA_X1_LVT frontend_0_i_124_12 (.CO(frontend_0_n_124_12), .S(
      frontend_0_pc_incr[13]), .A(pc[13]), .B(frontend_0_n_124_11));
  HA_X1_LVT frontend_0_i_124_13 (.CO(frontend_0_n_124_13), .S(
      frontend_0_pc_incr[14]), .A(pc[14]), .B(frontend_0_n_124_12));
  XNOR2_X1_LVT frontend_0_i_124_14 (.ZN(frontend_0_n_124_14), .A(pc[15]), .B(
      frontend_0_n_124_13));
  INV_X1_LVT frontend_0_i_124_15 (.ZN(frontend_0_pc_incr[15]), .A(
      frontend_0_n_124_14));
  AOI221_X1_LVT frontend_0_i_126_30 (.ZN(frontend_0_n_126_15), .A(
      frontend_0_n_221), .B1(frontend_0_n_220), .B2(fe_mdb_in[15]), .C1(
      frontend_0_n_222), .C2(frontend_0_pc_incr[15]));
  INV_X1_LVT frontend_0_i_126_31 (.ZN(frontend_0_n_238), .A(frontend_0_n_126_15));
  AOI22_X1_LVT frontend_0_i_127_31 (.ZN(frontend_0_n_127_16), .A1(
      frontend_0_n_127_0), .A2(frontend_0_n_238), .B1(pc_sw_wr), .B2(pc_sw[15]));
  INV_X1_LVT frontend_0_i_127_32 (.ZN(pc_nxt[15]), .A(frontend_0_n_127_16));
  DFFR_X1_LVT \frontend_0_pc_reg[0] (.Q(pc[0]), .QN(), .CK(cpu_mclk), .D(pc_nxt[0]), 
      .RN(frontend_0_n_91));
  AOI22_X1_LVT frontend_0_i_126_0 (.ZN(frontend_0_n_126_0), .A1(fe_mdb_in[0]), 
      .A2(frontend_0_n_220), .B1(pc[0]), .B2(frontend_0_n_222));
  INV_X1_LVT frontend_0_i_126_1 (.ZN(frontend_0_n_223), .A(frontend_0_n_126_0));
  AOI22_X1_LVT frontend_0_i_127_1 (.ZN(frontend_0_n_127_1), .A1(
      frontend_0_n_127_0), .A2(frontend_0_n_223), .B1(pc_sw[0]), .B2(pc_sw_wr));
  INV_X1_LVT frontend_0_i_127_2 (.ZN(pc_nxt[0]), .A(frontend_0_n_127_1));
  DFFR_X1_LVT frontend_0_pmem_busy_reg (.Q(frontend_0_pmem_busy), .QN(), .CK(
      cpu_mclk), .D(fe_pmem_wait), .RN(frontend_0_n_91));
  NOR4_X1_LVT frontend_0_i_128_0 (.ZN(frontend_0_n_128_0), .A1(pc_sw_wr), .A2(
      frontend_0_fetch), .A3(frontend_0_pmem_busy), .A4(frontend_0_n_8));
  NAND2_X1_LVT frontend_0_i_128_1 (.ZN(frontend_0_n_128_1), .A1(cpu_halt_st), 
      .A2(frontend_0_n_0));
  NAND2_X1_LVT frontend_0_i_128_2 (.ZN(fe_mb_en), .A1(frontend_0_n_128_0), .A2(
      frontend_0_n_128_1));
  AND2_X1_LVT frontend_0_i_129_0 (.ZN(mclk_dma_enable), .A1(dma_en), .A2(
      cpu_en_s));
  AND2_X1_LVT frontend_0_and_mclk_dma_wkup_i_0_0 (.ZN(mclk_dma_wkup), .A1(
      dma_wkup), .A2(cpu_en_s));
  INV_X1_LVT frontend_0_i_130_0 (.ZN(frontend_0_n_130_0), .A(cpu_en_s));
  OAI211_X1_LVT frontend_0_i_130_1 (.ZN(frontend_0_n_130_1), .A(frontend_0_n_5), 
      .B(frontend_0_n_67), .C1(frontend_0_n_130_0), .C2(cpuoff));
  INV_X1_LVT frontend_0_i_130_2 (.ZN(frontend_0_n_130_2), .A(inst_irq_rst));
  AOI22_X1_LVT frontend_0_i_130_3 (.ZN(frontend_0_n_130_3), .A1(
      frontend_0_n_130_1), .A2(frontend_0_n_130_2), .B1(cpu_en_s), .B2(
      inst_irq_rst));
  INV_X1_LVT frontend_0_i_130_4 (.ZN(mclk_enable), .A(frontend_0_n_130_3));
  OR2_X1_LVT frontend_0_i_132_0 (.ZN(frontend_0_n_240), .A1(wkup), .A2(wdt_wkup));
  AND2_X1_LVT frontend_0_and_mirq_wkup_i_0_0 (.ZN(frontend_0_mirq_wkup), .A1(
      frontend_0_n_240), .A2(gie));
  OR2_X1_LVT frontend_0_i_131_0 (.ZN(frontend_0_n_239), .A1(nmi_wkup), .A2(
      frontend_0_mirq_wkup));
  AND2_X1_LVT frontend_0_and_mclk_wkup_i_0_0 (.ZN(mclk_wkup), .A1(
      frontend_0_n_239), .A2(cpu_en_s));
  NOR2_X1_LVT frontend_0_i_120_35 (.ZN(frontend_0_n_219), .A1(
      frontend_0_n_120_13), .A2(frontend_0_n_120_20));
  AND2_X1_LVT frontend_0_i_121_14 (.ZN(nmi_acc), .A1(frontend_0_n_8), .A2(
      frontend_0_n_219));
  INV_X1_LVT execution_unit_0_i_0_0 (.ZN(execution_unit_0_n_0_0), .A(e_state[3]));
  INV_X1_LVT execution_unit_0_i_0_1 (.ZN(execution_unit_0_n_0_1), .A(e_state[0]));
  INV_X1_LVT execution_unit_0_i_0_2 (.ZN(execution_unit_0_n_0_2), .A(e_state[1]));
  NOR4_X1_LVT execution_unit_0_i_0_3 (.ZN(execution_unit_0_n_0), .A1(
      execution_unit_0_n_0_0), .A2(execution_unit_0_n_0_1), .A3(
      execution_unit_0_n_0_2), .A4(e_state[2]));
  OR3_X1_LVT execution_unit_0_i_38_0 (.ZN(execution_unit_0_n_69), .A1(inst_as[4]), 
      .A2(inst_as[1]), .A3(inst_as[6]));
  INV_X1_LVT execution_unit_0_i_0_4 (.ZN(execution_unit_0_n_0_3), .A(e_state[2]));
  NOR4_X1_LVT execution_unit_0_i_0_5 (.ZN(execution_unit_0_n_1), .A1(
      execution_unit_0_n_0_2), .A2(execution_unit_0_n_0_3), .A3(e_state[0]), .A4(
      e_state[3]));
  NOR4_X1_LVT execution_unit_0_i_0_6 (.ZN(execution_unit_0_n_2), .A1(
      execution_unit_0_n_0_3), .A2(execution_unit_0_n_0_1), .A3(
      execution_unit_0_n_0_2), .A4(e_state[3]));
  AOI22_X1_LVT execution_unit_0_i_39_11 (.ZN(execution_unit_0_n_39_8), .A1(
      execution_unit_0_n_69), .A2(execution_unit_0_n_1), .B1(
      execution_unit_0_n_69), .B2(execution_unit_0_n_2));
  INV_X1_LVT execution_unit_0_i_39_12 (.ZN(execution_unit_0_n_73), .A(
      execution_unit_0_n_39_8));
  INV_X1_LVT execution_unit_0_i_40_4 (.ZN(execution_unit_0_n_40_4), .A(
      execution_unit_0_n_73));
  NOR2_X1_LVT execution_unit_0_i_40_5 (.ZN(execution_unit_0_n_74), .A1(
      execution_unit_0_n_40_4), .A2(cpu_halt_st));
  NAND2_X1_LVT execution_unit_0_i_41_90 (.ZN(execution_unit_0_n_41_75), .A1(
      execution_unit_0_n_74), .A2(inst_sext[15]));
  OR2_X1_LVT execution_unit_0_i_40_0 (.ZN(execution_unit_0_n_40_0), .A1(
      execution_unit_0_n_73), .A2(cpu_halt_st));
  NOR4_X1_LVT execution_unit_0_i_0_7 (.ZN(execution_unit_0_n_3), .A1(
      execution_unit_0_n_0_2), .A2(execution_unit_0_n_0_0), .A3(e_state[0]), .A4(
      e_state[2]));
  AND2_X1_LVT execution_unit_0_i_22_0 (.ZN(execution_unit_0_n_40), .A1(
      inst_so[6]), .A2(execution_unit_0_n_3));
  INV_X1_LVT execution_unit_0_i_39_8 (.ZN(execution_unit_0_n_39_6), .A(
      execution_unit_0_n_40));
  INV_X1_LVT execution_unit_0_i_2_0 (.ZN(execution_unit_0_n_10), .A(inst_so[6]));
  AND2_X1_LVT execution_unit_0_i_36_0 (.ZN(execution_unit_0_n_67), .A1(
      execution_unit_0_n_0), .A2(execution_unit_0_n_10));
  INV_X1_LVT execution_unit_0_i_39_9 (.ZN(execution_unit_0_n_39_7), .A(
      execution_unit_0_n_67));
  OR3_X1_LVT execution_unit_0_i_37_0 (.ZN(execution_unit_0_n_68), .A1(inst_ad[0]), 
      .A2(inst_type[0]), .A3(inst_type[1]));
  OAI21_X1_LVT execution_unit_0_i_39_10 (.ZN(execution_unit_0_n_72), .A(
      execution_unit_0_n_39_6), .B1(execution_unit_0_n_39_7), .B2(
      execution_unit_0_n_68));
  INV_X1_LVT execution_unit_0_i_40_6 (.ZN(execution_unit_0_n_40_5), .A(
      execution_unit_0_n_72));
  NOR2_X1_LVT execution_unit_0_i_40_7 (.ZN(execution_unit_0_n_75), .A1(
      execution_unit_0_n_40_0), .A2(execution_unit_0_n_40_5));
  INV_X1_LVT execution_unit_0_i_33_0 (.ZN(execution_unit_0_n_47), .A(inst_bw));
  INV_X1_LVT execution_unit_0_i_6_0 (.ZN(execution_unit_0_n_13), .A(inst_alu[11]));
  INV_X1_LVT execution_unit_0_i_3_0 (.ZN(execution_unit_0_n_11), .A(inst_irq_rst));
  NOR4_X1_LVT execution_unit_0_i_0_10 (.ZN(execution_unit_0_n_6), .A1(
      execution_unit_0_n_0_1), .A2(execution_unit_0_n_0_2), .A3(e_state[2]), .A4(
      e_state[3]));
  NOR4_X1_LVT execution_unit_0_i_0_9 (.ZN(execution_unit_0_n_5), .A1(
      execution_unit_0_n_0_1), .A2(e_state[1]), .A3(e_state[2]), .A4(e_state[3]));
  OAI21_X1_LVT execution_unit_0_i_4_0 (.ZN(execution_unit_0_n_4_0), .A(
      execution_unit_0_n_11), .B1(execution_unit_0_n_6), .B2(
      execution_unit_0_n_5));
  NAND2_X1_LVT execution_unit_0_i_4_1 (.ZN(execution_unit_0_n_4_1), .A1(
      execution_unit_0_n_10), .A2(execution_unit_0_n_3));
  NAND2_X1_LVT execution_unit_0_i_4_2 (.ZN(execution_unit_0_n_12), .A1(
      execution_unit_0_n_4_0), .A2(execution_unit_0_n_4_1));
  OR2_X1_LVT execution_unit_0_i_5_0 (.ZN(execution_unit_0_mb_wr_det), .A1(
      execution_unit_0_n_12), .A2(execution_unit_0_n_2));
  AND2_X1_LVT execution_unit_0_i_7_0 (.ZN(execution_unit_0_n_7_0), .A1(
      execution_unit_0_n_13), .A2(execution_unit_0_mb_wr_det));
  NOR4_X1_LVT execution_unit_0_i_0_8 (.ZN(execution_unit_0_n_4), .A1(
      execution_unit_0_n_0_1), .A2(execution_unit_0_n_0_0), .A3(e_state[1]), .A4(
      e_state[2]));
  INV_X1_LVT execution_unit_0_i_7_1 (.ZN(execution_unit_0_n_7_1), .A(
      execution_unit_0_n_4));
  NOR3_X1_LVT execution_unit_0_i_7_2 (.ZN(execution_unit_0_n_7_2), .A1(
      execution_unit_0_n_7_1), .A2(inst_type[0]), .A3(inst_mov));
  INV_X1_LVT execution_unit_0_i_7_3 (.ZN(execution_unit_0_n_7_3), .A(
      execution_unit_0_n_1));
  NOR2_X1_LVT execution_unit_0_i_7_4 (.ZN(execution_unit_0_n_7_4), .A1(
      execution_unit_0_n_7_3), .A2(inst_as[5]));
  AND2_X1_LVT execution_unit_0_i_1_0 (.ZN(execution_unit_0_n_9), .A1(
      execution_unit_0_n_0), .A2(inst_so[6]));
  OR4_X1_LVT execution_unit_0_i_7_5 (.ZN(eu_mb_en), .A1(execution_unit_0_n_7_0), 
      .A2(execution_unit_0_n_7_2), .A3(execution_unit_0_n_7_4), .A4(
      execution_unit_0_n_9));
  CLKGATETST_X1_LVT execution_unit_0_clk_gate_mab_lsb_reg (.GCK(
      execution_unit_0_n_16), .CK(cpu_mclk), .E(eu_mb_en), .SE(1'b0));
  INV_X1_LVT execution_unit_0_i_11_0 (.ZN(execution_unit_0_n_18), .A(puc_rst));
  DFFR_X1_LVT execution_unit_0_mab_lsb_reg (.Q(execution_unit_0_mab_lsb), .QN(), 
      .CK(execution_unit_0_n_16), .D(eu_mab[0]), .RN(execution_unit_0_n_18));
  AND2_X1_LVT execution_unit_0_i_33_2 (.ZN(execution_unit_0_n_49), .A1(
      execution_unit_0_mab_lsb), .A2(inst_bw));
  NOR2_X1_LVT execution_unit_0_i_33_1 (.ZN(execution_unit_0_n_48), .A1(
      execution_unit_0_n_47), .A2(execution_unit_0_mab_lsb));
  NOR3_X1_LVT execution_unit_0_i_34_17 (.ZN(execution_unit_0_n_34_9), .A1(
      execution_unit_0_n_47), .A2(execution_unit_0_n_49), .A3(
      execution_unit_0_n_48));
  INV_X1_LVT execution_unit_0_i_34_32 (.ZN(execution_unit_0_n_34_17), .A(
      eu_mdb_in[15]));
  NOR2_X1_LVT execution_unit_0_i_34_33 (.ZN(execution_unit_0_n_65), .A1(
      execution_unit_0_n_34_9), .A2(execution_unit_0_n_34_17));
  NAND2_X1_LVT execution_unit_0_i_41_91 (.ZN(execution_unit_0_n_41_76), .A1(
      execution_unit_0_n_75), .A2(execution_unit_0_n_65));
  NOR2_X1_LVT execution_unit_0_i_40_1 (.ZN(execution_unit_0_n_40_1), .A1(
      execution_unit_0_n_40_0), .A2(execution_unit_0_n_72));
  INV_X1_LVT execution_unit_0_i_39_3 (.ZN(execution_unit_0_n_39_2), .A(
      execution_unit_0_n_4));
  OR2_X1_LVT execution_unit_0_i_18_0 (.ZN(execution_unit_0_n_37), .A1(inst_so[4]), 
      .A2(inst_so[5]));
  OR2_X1_LVT execution_unit_0_i_19_0 (.ZN(execution_unit_0_n_38), .A1(inst_so[6]), 
      .A2(execution_unit_0_n_37));
  NOR3_X1_LVT execution_unit_0_i_39_4 (.ZN(execution_unit_0_n_39_3), .A1(
      execution_unit_0_n_39_2), .A2(inst_ad[6]), .A3(execution_unit_0_n_38));
  INV_X1_LVT execution_unit_0_i_39_5 (.ZN(execution_unit_0_n_39_4), .A(
      inst_ad[6]));
  AOI221_X1_LVT execution_unit_0_i_39_6 (.ZN(execution_unit_0_n_39_5), .A(
      execution_unit_0_n_39_3), .B1(execution_unit_0_n_39_4), .B2(
      execution_unit_0_n_3), .C1(execution_unit_0_n_68), .C2(
      execution_unit_0_n_67));
  INV_X1_LVT execution_unit_0_i_39_7 (.ZN(execution_unit_0_n_71), .A(
      execution_unit_0_n_39_5));
  AND2_X1_LVT execution_unit_0_i_40_8 (.ZN(execution_unit_0_n_76), .A1(
      execution_unit_0_n_40_1), .A2(execution_unit_0_n_71));
  NAND2_X1_LVT execution_unit_0_i_41_92 (.ZN(execution_unit_0_n_41_77), .A1(
      execution_unit_0_n_76), .A2(dbg_reg_din[15]));
  INV_X1_LVT execution_unit_0_i_40_2 (.ZN(execution_unit_0_n_40_2), .A(
      execution_unit_0_n_71));
  NAND2_X1_LVT execution_unit_0_i_40_3 (.ZN(execution_unit_0_n_40_3), .A1(
      execution_unit_0_n_40_1), .A2(execution_unit_0_n_40_2));
  OR2_X1_LVT execution_unit_0_i_24_0 (.ZN(execution_unit_0_n_41), .A1(inst_as[2]), 
      .A2(inst_as[3]));
  AND2_X1_LVT execution_unit_0_i_25_0 (.ZN(execution_unit_0_n_42), .A1(
      inst_src[1]), .A2(execution_unit_0_n_41));
  AND3_X1_LVT execution_unit_0_i_26_0 (.ZN(execution_unit_0_n_43), .A1(
      execution_unit_0_n_42), .A2(execution_unit_0_n_1), .A3(
      execution_unit_0_n_37));
  NOR4_X1_LVT execution_unit_0_i_0_12 (.ZN(execution_unit_0_n_8), .A1(
      execution_unit_0_n_0_1), .A2(execution_unit_0_n_0_3), .A3(e_state[1]), .A4(
      e_state[3]));
  AND3_X1_LVT execution_unit_0_i_27_0 (.ZN(execution_unit_0_n_44), .A1(
      inst_as[1]), .A2(execution_unit_0_n_8), .A3(execution_unit_0_n_37));
  OR2_X1_LVT execution_unit_0_i_29_0 (.ZN(execution_unit_0_n_46), .A1(
      execution_unit_0_n_5), .A2(execution_unit_0_n_6));
  OR2_X1_LVT execution_unit_0_i_35_0 (.ZN(execution_unit_0_n_66), .A1(
      execution_unit_0_n_44), .A2(execution_unit_0_n_46));
  NOR4_X1_LVT execution_unit_0_i_0_11 (.ZN(execution_unit_0_n_7), .A1(
      execution_unit_0_n_0_2), .A2(e_state[0]), .A3(e_state[2]), .A4(e_state[3]));
  NOR3_X1_LVT execution_unit_0_i_39_0 (.ZN(execution_unit_0_n_39_0), .A1(
      execution_unit_0_n_43), .A2(execution_unit_0_n_66), .A3(
      execution_unit_0_n_7));
  AND2_X1_LVT execution_unit_0_i_28_0 (.ZN(execution_unit_0_n_45), .A1(
      execution_unit_0_n_37), .A2(execution_unit_0_n_4));
  NAND2_X1_LVT execution_unit_0_i_39_1 (.ZN(execution_unit_0_n_39_1), .A1(
      execution_unit_0_n_10), .A2(execution_unit_0_n_45));
  NAND2_X1_LVT execution_unit_0_i_39_2 (.ZN(execution_unit_0_n_70), .A1(
      execution_unit_0_n_39_0), .A2(execution_unit_0_n_39_1));
  INV_X1_LVT execution_unit_0_i_40_9 (.ZN(execution_unit_0_n_40_6), .A(
      execution_unit_0_n_70));
  NOR2_X1_LVT execution_unit_0_i_40_10 (.ZN(execution_unit_0_n_77), .A1(
      execution_unit_0_n_40_3), .A2(execution_unit_0_n_40_6));
  INV_X1_LVT execution_unit_0_i_41_8 (.ZN(execution_unit_0_n_41_7), .A(
      execution_unit_0_n_77));
  NAND4_X1_LVT execution_unit_0_i_41_93 (.ZN(execution_unit_0_n_41_78), .A1(
      execution_unit_0_n_41_75), .A2(execution_unit_0_n_41_76), .A3(
      execution_unit_0_n_41_77), .A4(execution_unit_0_n_41_7));
  AOI21_X1_LVT execution_unit_0_i_41_94 (.ZN(execution_unit_0_n_41_79), .A(
      execution_unit_0_n_41_78), .B1(cpu_halt_st), .B2(dbg_mem_dout[15]));
  INV_X1_LVT execution_unit_0_i_41_95 (.ZN(execution_unit_0_n_93), .A(
      execution_unit_0_n_41_79));
  NAND2_X1_LVT execution_unit_0_i_41_84 (.ZN(execution_unit_0_n_41_70), .A1(
      execution_unit_0_n_74), .A2(inst_sext[14]));
  INV_X1_LVT execution_unit_0_i_34_30 (.ZN(execution_unit_0_n_34_16), .A(
      eu_mdb_in[14]));
  NOR2_X1_LVT execution_unit_0_i_34_31 (.ZN(execution_unit_0_n_64), .A1(
      execution_unit_0_n_34_9), .A2(execution_unit_0_n_34_16));
  NAND2_X1_LVT execution_unit_0_i_41_85 (.ZN(execution_unit_0_n_41_71), .A1(
      execution_unit_0_n_75), .A2(execution_unit_0_n_64));
  NAND2_X1_LVT execution_unit_0_i_41_86 (.ZN(execution_unit_0_n_41_72), .A1(
      execution_unit_0_n_76), .A2(dbg_reg_din[14]));
  NAND4_X1_LVT execution_unit_0_i_41_87 (.ZN(execution_unit_0_n_41_73), .A1(
      execution_unit_0_n_41_70), .A2(execution_unit_0_n_41_71), .A3(
      execution_unit_0_n_41_72), .A4(execution_unit_0_n_41_7));
  AOI21_X1_LVT execution_unit_0_i_41_88 (.ZN(execution_unit_0_n_41_74), .A(
      execution_unit_0_n_41_73), .B1(cpu_halt_st), .B2(dbg_mem_dout[14]));
  INV_X1_LVT execution_unit_0_i_41_89 (.ZN(execution_unit_0_n_92), .A(
      execution_unit_0_n_41_74));
  NAND2_X1_LVT execution_unit_0_i_41_78 (.ZN(execution_unit_0_n_41_65), .A1(
      execution_unit_0_n_74), .A2(inst_sext[13]));
  INV_X1_LVT execution_unit_0_i_34_28 (.ZN(execution_unit_0_n_34_15), .A(
      eu_mdb_in[13]));
  NOR2_X1_LVT execution_unit_0_i_34_29 (.ZN(execution_unit_0_n_63), .A1(
      execution_unit_0_n_34_9), .A2(execution_unit_0_n_34_15));
  NAND2_X1_LVT execution_unit_0_i_41_79 (.ZN(execution_unit_0_n_41_66), .A1(
      execution_unit_0_n_75), .A2(execution_unit_0_n_63));
  NAND2_X1_LVT execution_unit_0_i_41_80 (.ZN(execution_unit_0_n_41_67), .A1(
      execution_unit_0_n_76), .A2(dbg_reg_din[13]));
  NAND4_X1_LVT execution_unit_0_i_41_81 (.ZN(execution_unit_0_n_41_68), .A1(
      execution_unit_0_n_41_65), .A2(execution_unit_0_n_41_66), .A3(
      execution_unit_0_n_41_67), .A4(execution_unit_0_n_41_7));
  AOI21_X1_LVT execution_unit_0_i_41_82 (.ZN(execution_unit_0_n_41_69), .A(
      execution_unit_0_n_41_68), .B1(cpu_halt_st), .B2(dbg_mem_dout[13]));
  INV_X1_LVT execution_unit_0_i_41_83 (.ZN(execution_unit_0_n_91), .A(
      execution_unit_0_n_41_69));
  NAND2_X1_LVT execution_unit_0_i_41_72 (.ZN(execution_unit_0_n_41_60), .A1(
      execution_unit_0_n_74), .A2(inst_sext[12]));
  INV_X1_LVT execution_unit_0_i_34_26 (.ZN(execution_unit_0_n_34_14), .A(
      eu_mdb_in[12]));
  NOR2_X1_LVT execution_unit_0_i_34_27 (.ZN(execution_unit_0_n_62), .A1(
      execution_unit_0_n_34_9), .A2(execution_unit_0_n_34_14));
  NAND2_X1_LVT execution_unit_0_i_41_73 (.ZN(execution_unit_0_n_41_61), .A1(
      execution_unit_0_n_75), .A2(execution_unit_0_n_62));
  NAND2_X1_LVT execution_unit_0_i_41_74 (.ZN(execution_unit_0_n_41_62), .A1(
      execution_unit_0_n_76), .A2(dbg_reg_din[12]));
  NAND4_X1_LVT execution_unit_0_i_41_75 (.ZN(execution_unit_0_n_41_63), .A1(
      execution_unit_0_n_41_60), .A2(execution_unit_0_n_41_61), .A3(
      execution_unit_0_n_41_62), .A4(execution_unit_0_n_41_7));
  AOI21_X1_LVT execution_unit_0_i_41_76 (.ZN(execution_unit_0_n_41_64), .A(
      execution_unit_0_n_41_63), .B1(cpu_halt_st), .B2(dbg_mem_dout[12]));
  INV_X1_LVT execution_unit_0_i_41_77 (.ZN(execution_unit_0_n_90), .A(
      execution_unit_0_n_41_64));
  NAND2_X1_LVT execution_unit_0_i_41_66 (.ZN(execution_unit_0_n_41_55), .A1(
      execution_unit_0_n_74), .A2(inst_sext[11]));
  INV_X1_LVT execution_unit_0_i_34_24 (.ZN(execution_unit_0_n_34_13), .A(
      eu_mdb_in[11]));
  NOR2_X1_LVT execution_unit_0_i_34_25 (.ZN(execution_unit_0_n_61), .A1(
      execution_unit_0_n_34_9), .A2(execution_unit_0_n_34_13));
  NAND2_X1_LVT execution_unit_0_i_41_67 (.ZN(execution_unit_0_n_41_56), .A1(
      execution_unit_0_n_75), .A2(execution_unit_0_n_61));
  NAND2_X1_LVT execution_unit_0_i_41_68 (.ZN(execution_unit_0_n_41_57), .A1(
      execution_unit_0_n_76), .A2(dbg_reg_din[11]));
  NAND4_X1_LVT execution_unit_0_i_41_69 (.ZN(execution_unit_0_n_41_58), .A1(
      execution_unit_0_n_41_55), .A2(execution_unit_0_n_41_56), .A3(
      execution_unit_0_n_41_57), .A4(execution_unit_0_n_41_7));
  AOI21_X1_LVT execution_unit_0_i_41_70 (.ZN(execution_unit_0_n_41_59), .A(
      execution_unit_0_n_41_58), .B1(cpu_halt_st), .B2(dbg_mem_dout[11]));
  INV_X1_LVT execution_unit_0_i_41_71 (.ZN(execution_unit_0_n_89), .A(
      execution_unit_0_n_41_59));
  NAND2_X1_LVT execution_unit_0_i_41_60 (.ZN(execution_unit_0_n_41_50), .A1(
      execution_unit_0_n_74), .A2(inst_sext[10]));
  INV_X1_LVT execution_unit_0_i_34_22 (.ZN(execution_unit_0_n_34_12), .A(
      eu_mdb_in[10]));
  NOR2_X1_LVT execution_unit_0_i_34_23 (.ZN(execution_unit_0_n_60), .A1(
      execution_unit_0_n_34_9), .A2(execution_unit_0_n_34_12));
  NAND2_X1_LVT execution_unit_0_i_41_61 (.ZN(execution_unit_0_n_41_51), .A1(
      execution_unit_0_n_75), .A2(execution_unit_0_n_60));
  NAND2_X1_LVT execution_unit_0_i_41_62 (.ZN(execution_unit_0_n_41_52), .A1(
      execution_unit_0_n_76), .A2(dbg_reg_din[10]));
  NAND4_X1_LVT execution_unit_0_i_41_63 (.ZN(execution_unit_0_n_41_53), .A1(
      execution_unit_0_n_41_50), .A2(execution_unit_0_n_41_51), .A3(
      execution_unit_0_n_41_52), .A4(execution_unit_0_n_41_7));
  AOI21_X1_LVT execution_unit_0_i_41_64 (.ZN(execution_unit_0_n_41_54), .A(
      execution_unit_0_n_41_53), .B1(cpu_halt_st), .B2(dbg_mem_dout[10]));
  INV_X1_LVT execution_unit_0_i_41_65 (.ZN(execution_unit_0_n_88), .A(
      execution_unit_0_n_41_54));
  NAND2_X1_LVT execution_unit_0_i_41_54 (.ZN(execution_unit_0_n_41_45), .A1(
      execution_unit_0_n_74), .A2(inst_sext[9]));
  INV_X1_LVT execution_unit_0_i_34_20 (.ZN(execution_unit_0_n_34_11), .A(
      eu_mdb_in[9]));
  NOR2_X1_LVT execution_unit_0_i_34_21 (.ZN(execution_unit_0_n_59), .A1(
      execution_unit_0_n_34_9), .A2(execution_unit_0_n_34_11));
  NAND2_X1_LVT execution_unit_0_i_41_55 (.ZN(execution_unit_0_n_41_46), .A1(
      execution_unit_0_n_75), .A2(execution_unit_0_n_59));
  NAND2_X1_LVT execution_unit_0_i_41_56 (.ZN(execution_unit_0_n_41_47), .A1(
      execution_unit_0_n_76), .A2(dbg_reg_din[9]));
  NAND4_X1_LVT execution_unit_0_i_41_57 (.ZN(execution_unit_0_n_41_48), .A1(
      execution_unit_0_n_41_45), .A2(execution_unit_0_n_41_46), .A3(
      execution_unit_0_n_41_47), .A4(execution_unit_0_n_41_7));
  AOI21_X1_LVT execution_unit_0_i_41_58 (.ZN(execution_unit_0_n_41_49), .A(
      execution_unit_0_n_41_48), .B1(cpu_halt_st), .B2(dbg_mem_dout[9]));
  INV_X1_LVT execution_unit_0_i_41_59 (.ZN(execution_unit_0_n_87), .A(
      execution_unit_0_n_41_49));
  NAND2_X1_LVT execution_unit_0_i_41_48 (.ZN(execution_unit_0_n_41_40), .A1(
      execution_unit_0_n_74), .A2(inst_sext[8]));
  INV_X1_LVT execution_unit_0_i_34_18 (.ZN(execution_unit_0_n_34_10), .A(
      eu_mdb_in[8]));
  NOR2_X1_LVT execution_unit_0_i_34_19 (.ZN(execution_unit_0_n_58), .A1(
      execution_unit_0_n_34_9), .A2(execution_unit_0_n_34_10));
  NAND2_X1_LVT execution_unit_0_i_41_49 (.ZN(execution_unit_0_n_41_41), .A1(
      execution_unit_0_n_75), .A2(execution_unit_0_n_58));
  NAND2_X1_LVT execution_unit_0_i_41_50 (.ZN(execution_unit_0_n_41_42), .A1(
      execution_unit_0_n_76), .A2(dbg_reg_din[8]));
  NAND4_X1_LVT execution_unit_0_i_41_51 (.ZN(execution_unit_0_n_41_43), .A1(
      execution_unit_0_n_41_40), .A2(execution_unit_0_n_41_41), .A3(
      execution_unit_0_n_41_42), .A4(execution_unit_0_n_41_7));
  AOI21_X1_LVT execution_unit_0_i_41_52 (.ZN(execution_unit_0_n_41_44), .A(
      execution_unit_0_n_41_43), .B1(cpu_halt_st), .B2(dbg_mem_dout[8]));
  INV_X1_LVT execution_unit_0_i_41_53 (.ZN(execution_unit_0_n_86), .A(
      execution_unit_0_n_41_44));
  NAND2_X1_LVT execution_unit_0_i_41_42 (.ZN(execution_unit_0_n_41_35), .A1(
      execution_unit_0_n_74), .A2(inst_sext[7]));
  OR2_X1_LVT execution_unit_0_i_34_0 (.ZN(execution_unit_0_n_34_0), .A1(
      execution_unit_0_n_47), .A2(execution_unit_0_n_48));
  AOI22_X1_LVT execution_unit_0_i_34_15 (.ZN(execution_unit_0_n_34_8), .A1(
      execution_unit_0_n_34_0), .A2(eu_mdb_in[7]), .B1(execution_unit_0_n_49), 
      .B2(eu_mdb_in[15]));
  INV_X1_LVT execution_unit_0_i_34_16 (.ZN(execution_unit_0_n_57), .A(
      execution_unit_0_n_34_8));
  NAND2_X1_LVT execution_unit_0_i_41_43 (.ZN(execution_unit_0_n_41_36), .A1(
      execution_unit_0_n_75), .A2(execution_unit_0_n_57));
  NAND2_X1_LVT execution_unit_0_i_41_44 (.ZN(execution_unit_0_n_41_37), .A1(
      execution_unit_0_n_76), .A2(dbg_reg_din[7]));
  NAND4_X1_LVT execution_unit_0_i_41_45 (.ZN(execution_unit_0_n_41_38), .A1(
      execution_unit_0_n_41_35), .A2(execution_unit_0_n_41_36), .A3(
      execution_unit_0_n_41_37), .A4(execution_unit_0_n_41_7));
  AOI21_X1_LVT execution_unit_0_i_41_46 (.ZN(execution_unit_0_n_41_39), .A(
      execution_unit_0_n_41_38), .B1(cpu_halt_st), .B2(dbg_mem_dout[7]));
  INV_X1_LVT execution_unit_0_i_41_47 (.ZN(execution_unit_0_n_85), .A(
      execution_unit_0_n_41_39));
  NAND2_X1_LVT execution_unit_0_i_41_36 (.ZN(execution_unit_0_n_41_30), .A1(
      execution_unit_0_n_74), .A2(inst_sext[6]));
  AOI22_X1_LVT execution_unit_0_i_34_13 (.ZN(execution_unit_0_n_34_7), .A1(
      execution_unit_0_n_34_0), .A2(eu_mdb_in[6]), .B1(execution_unit_0_n_49), 
      .B2(eu_mdb_in[14]));
  INV_X1_LVT execution_unit_0_i_34_14 (.ZN(execution_unit_0_n_56), .A(
      execution_unit_0_n_34_7));
  NAND2_X1_LVT execution_unit_0_i_41_37 (.ZN(execution_unit_0_n_41_31), .A1(
      execution_unit_0_n_75), .A2(execution_unit_0_n_56));
  NAND2_X1_LVT execution_unit_0_i_41_38 (.ZN(execution_unit_0_n_41_32), .A1(
      execution_unit_0_n_76), .A2(dbg_reg_din[6]));
  NAND4_X1_LVT execution_unit_0_i_41_39 (.ZN(execution_unit_0_n_41_33), .A1(
      execution_unit_0_n_41_30), .A2(execution_unit_0_n_41_31), .A3(
      execution_unit_0_n_41_32), .A4(execution_unit_0_n_41_7));
  AOI21_X1_LVT execution_unit_0_i_41_40 (.ZN(execution_unit_0_n_41_34), .A(
      execution_unit_0_n_41_33), .B1(cpu_halt_st), .B2(dbg_mem_dout[6]));
  INV_X1_LVT execution_unit_0_i_41_41 (.ZN(execution_unit_0_n_84), .A(
      execution_unit_0_n_41_34));
  NAND2_X1_LVT execution_unit_0_i_41_30 (.ZN(execution_unit_0_n_41_25), .A1(
      execution_unit_0_n_74), .A2(inst_sext[5]));
  AOI22_X1_LVT execution_unit_0_i_34_11 (.ZN(execution_unit_0_n_34_6), .A1(
      execution_unit_0_n_34_0), .A2(eu_mdb_in[5]), .B1(execution_unit_0_n_49), 
      .B2(eu_mdb_in[13]));
  INV_X1_LVT execution_unit_0_i_34_12 (.ZN(execution_unit_0_n_55), .A(
      execution_unit_0_n_34_6));
  NAND2_X1_LVT execution_unit_0_i_41_31 (.ZN(execution_unit_0_n_41_26), .A1(
      execution_unit_0_n_75), .A2(execution_unit_0_n_55));
  NAND2_X1_LVT execution_unit_0_i_41_32 (.ZN(execution_unit_0_n_41_27), .A1(
      execution_unit_0_n_76), .A2(dbg_reg_din[5]));
  NAND4_X1_LVT execution_unit_0_i_41_33 (.ZN(execution_unit_0_n_41_28), .A1(
      execution_unit_0_n_41_25), .A2(execution_unit_0_n_41_26), .A3(
      execution_unit_0_n_41_27), .A4(execution_unit_0_n_41_7));
  AOI21_X1_LVT execution_unit_0_i_41_34 (.ZN(execution_unit_0_n_41_29), .A(
      execution_unit_0_n_41_28), .B1(cpu_halt_st), .B2(dbg_mem_dout[5]));
  INV_X1_LVT execution_unit_0_i_41_35 (.ZN(execution_unit_0_n_83), .A(
      execution_unit_0_n_41_29));
  NAND2_X1_LVT execution_unit_0_i_41_24 (.ZN(execution_unit_0_n_41_20), .A1(
      execution_unit_0_n_74), .A2(inst_sext[4]));
  AOI22_X1_LVT execution_unit_0_i_34_9 (.ZN(execution_unit_0_n_34_5), .A1(
      execution_unit_0_n_34_0), .A2(eu_mdb_in[4]), .B1(execution_unit_0_n_49), 
      .B2(eu_mdb_in[12]));
  INV_X1_LVT execution_unit_0_i_34_10 (.ZN(execution_unit_0_n_54), .A(
      execution_unit_0_n_34_5));
  NAND2_X1_LVT execution_unit_0_i_41_25 (.ZN(execution_unit_0_n_41_21), .A1(
      execution_unit_0_n_75), .A2(execution_unit_0_n_54));
  NAND2_X1_LVT execution_unit_0_i_41_26 (.ZN(execution_unit_0_n_41_22), .A1(
      execution_unit_0_n_76), .A2(dbg_reg_din[4]));
  NAND4_X1_LVT execution_unit_0_i_41_27 (.ZN(execution_unit_0_n_41_23), .A1(
      execution_unit_0_n_41_20), .A2(execution_unit_0_n_41_21), .A3(
      execution_unit_0_n_41_22), .A4(execution_unit_0_n_41_7));
  AOI21_X1_LVT execution_unit_0_i_41_28 (.ZN(execution_unit_0_n_41_24), .A(
      execution_unit_0_n_41_23), .B1(cpu_halt_st), .B2(dbg_mem_dout[4]));
  INV_X1_LVT execution_unit_0_i_41_29 (.ZN(execution_unit_0_n_82), .A(
      execution_unit_0_n_41_24));
  NAND2_X1_LVT execution_unit_0_i_41_18 (.ZN(execution_unit_0_n_41_15), .A1(
      execution_unit_0_n_74), .A2(inst_sext[3]));
  AOI22_X1_LVT execution_unit_0_i_34_7 (.ZN(execution_unit_0_n_34_4), .A1(
      execution_unit_0_n_34_0), .A2(eu_mdb_in[3]), .B1(execution_unit_0_n_49), 
      .B2(eu_mdb_in[11]));
  INV_X1_LVT execution_unit_0_i_34_8 (.ZN(execution_unit_0_n_53), .A(
      execution_unit_0_n_34_4));
  NAND2_X1_LVT execution_unit_0_i_41_19 (.ZN(execution_unit_0_n_41_16), .A1(
      execution_unit_0_n_75), .A2(execution_unit_0_n_53));
  NAND2_X1_LVT execution_unit_0_i_41_20 (.ZN(execution_unit_0_n_41_17), .A1(
      execution_unit_0_n_76), .A2(dbg_reg_din[3]));
  NAND4_X1_LVT execution_unit_0_i_41_21 (.ZN(execution_unit_0_n_41_18), .A1(
      execution_unit_0_n_41_15), .A2(execution_unit_0_n_41_16), .A3(
      execution_unit_0_n_41_17), .A4(execution_unit_0_n_41_7));
  AOI21_X1_LVT execution_unit_0_i_41_22 (.ZN(execution_unit_0_n_41_19), .A(
      execution_unit_0_n_41_18), .B1(cpu_halt_st), .B2(dbg_mem_dout[3]));
  INV_X1_LVT execution_unit_0_i_41_23 (.ZN(execution_unit_0_n_81), .A(
      execution_unit_0_n_41_19));
  NAND2_X1_LVT execution_unit_0_i_41_12 (.ZN(execution_unit_0_n_41_10), .A1(
      execution_unit_0_n_74), .A2(inst_sext[2]));
  AOI22_X1_LVT execution_unit_0_i_34_5 (.ZN(execution_unit_0_n_34_3), .A1(
      execution_unit_0_n_34_0), .A2(eu_mdb_in[2]), .B1(execution_unit_0_n_49), 
      .B2(eu_mdb_in[10]));
  INV_X1_LVT execution_unit_0_i_34_6 (.ZN(execution_unit_0_n_52), .A(
      execution_unit_0_n_34_3));
  NAND2_X1_LVT execution_unit_0_i_41_13 (.ZN(execution_unit_0_n_41_11), .A1(
      execution_unit_0_n_75), .A2(execution_unit_0_n_52));
  NAND2_X1_LVT execution_unit_0_i_41_14 (.ZN(execution_unit_0_n_41_12), .A1(
      execution_unit_0_n_76), .A2(dbg_reg_din[2]));
  NAND4_X1_LVT execution_unit_0_i_41_15 (.ZN(execution_unit_0_n_41_13), .A1(
      execution_unit_0_n_41_10), .A2(execution_unit_0_n_41_11), .A3(
      execution_unit_0_n_41_12), .A4(execution_unit_0_n_41_7));
  AOI21_X1_LVT execution_unit_0_i_41_16 (.ZN(execution_unit_0_n_41_14), .A(
      execution_unit_0_n_41_13), .B1(cpu_halt_st), .B2(dbg_mem_dout[2]));
  INV_X1_LVT execution_unit_0_i_41_17 (.ZN(execution_unit_0_n_80), .A(
      execution_unit_0_n_41_14));
  NAND2_X1_LVT execution_unit_0_i_41_5 (.ZN(execution_unit_0_n_41_4), .A1(
      execution_unit_0_n_74), .A2(inst_sext[1]));
  AOI22_X1_LVT execution_unit_0_i_34_3 (.ZN(execution_unit_0_n_34_2), .A1(
      execution_unit_0_n_34_0), .A2(eu_mdb_in[1]), .B1(execution_unit_0_n_49), 
      .B2(eu_mdb_in[9]));
  INV_X1_LVT execution_unit_0_i_34_4 (.ZN(execution_unit_0_n_51), .A(
      execution_unit_0_n_34_2));
  NAND2_X1_LVT execution_unit_0_i_41_6 (.ZN(execution_unit_0_n_41_5), .A1(
      execution_unit_0_n_75), .A2(execution_unit_0_n_51));
  NAND2_X1_LVT execution_unit_0_i_41_7 (.ZN(execution_unit_0_n_41_6), .A1(
      execution_unit_0_n_76), .A2(dbg_reg_din[1]));
  NAND4_X1_LVT execution_unit_0_i_41_9 (.ZN(execution_unit_0_n_41_8), .A1(
      execution_unit_0_n_41_4), .A2(execution_unit_0_n_41_5), .A3(
      execution_unit_0_n_41_6), .A4(execution_unit_0_n_41_7));
  AOI21_X1_LVT execution_unit_0_i_41_10 (.ZN(execution_unit_0_n_41_9), .A(
      execution_unit_0_n_41_8), .B1(cpu_halt_st), .B2(dbg_mem_dout[1]));
  INV_X1_LVT execution_unit_0_i_41_11 (.ZN(execution_unit_0_n_79), .A(
      execution_unit_0_n_41_9));
  NAND2_X1_LVT execution_unit_0_i_41_0 (.ZN(execution_unit_0_n_41_0), .A1(
      dbg_mem_dout[0]), .A2(cpu_halt_st));
  NAND2_X1_LVT execution_unit_0_i_41_1 (.ZN(execution_unit_0_n_41_1), .A1(
      inst_sext[0]), .A2(execution_unit_0_n_74));
  AOI22_X1_LVT execution_unit_0_i_34_1 (.ZN(execution_unit_0_n_34_1), .A1(
      execution_unit_0_n_34_0), .A2(eu_mdb_in[0]), .B1(eu_mdb_in[8]), .B2(
      execution_unit_0_n_49));
  INV_X1_LVT execution_unit_0_i_34_2 (.ZN(execution_unit_0_n_50), .A(
      execution_unit_0_n_34_1));
  NAND2_X1_LVT execution_unit_0_i_41_2 (.ZN(execution_unit_0_n_41_2), .A1(
      execution_unit_0_n_50), .A2(execution_unit_0_n_75));
  NAND2_X1_LVT execution_unit_0_i_41_3 (.ZN(execution_unit_0_n_41_3), .A1(
      dbg_reg_din[0]), .A2(execution_unit_0_n_76));
  NAND4_X1_LVT execution_unit_0_i_41_4 (.ZN(execution_unit_0_n_78), .A1(
      execution_unit_0_n_41_0), .A2(execution_unit_0_n_41_1), .A3(
      execution_unit_0_n_41_2), .A4(execution_unit_0_n_41_3));
  OR2_X1_LVT execution_unit_0_i_48_8 (.ZN(execution_unit_0_n_102), .A1(
      execution_unit_0_n_45), .A2(execution_unit_0_n_66));
  NOR4_X1_LVT execution_unit_0_i_0_13 (.ZN(execution_unit_0_reg_sr_clr), .A1(
      e_state[0]), .A2(e_state[1]), .A3(e_state[2]), .A4(e_state[3]));
  NOR2_X1_LVT execution_unit_0_i_48_9 (.ZN(execution_unit_0_n_48_5), .A1(
      execution_unit_0_reg_sr_clr), .A2(execution_unit_0_n_7));
  INV_X1_LVT execution_unit_0_i_48_10 (.ZN(execution_unit_0_n_48_6), .A(
      inst_type[1]));
  NAND3_X1_LVT execution_unit_0_i_48_11 (.ZN(execution_unit_0_n_48_7), .A1(
      execution_unit_0_n_48_6), .A2(inst_as[0]), .A3(execution_unit_0_n_0));
  INV_X1_LVT execution_unit_0_i_47_0 (.ZN(execution_unit_0_n_98), .A(inst_as[6]));
  NAND2_X1_LVT execution_unit_0_i_48_12 (.ZN(execution_unit_0_n_48_8), .A1(
      execution_unit_0_n_2), .A2(execution_unit_0_n_98));
  NAND2_X1_LVT execution_unit_0_i_48_13 (.ZN(execution_unit_0_n_48_9), .A1(
      execution_unit_0_n_98), .A2(execution_unit_0_n_1));
  NAND4_X1_LVT execution_unit_0_i_48_14 (.ZN(execution_unit_0_n_103), .A1(
      execution_unit_0_n_48_5), .A2(execution_unit_0_n_48_7), .A3(
      execution_unit_0_n_48_8), .A4(execution_unit_0_n_48_9));
  NOR2_X1_LVT execution_unit_0_i_49_0 (.ZN(execution_unit_0_n_49_0), .A1(
      execution_unit_0_n_102), .A2(execution_unit_0_n_103));
  INV_X1_LVT execution_unit_0_i_49_8 (.ZN(execution_unit_0_n_49_7), .A(
      execution_unit_0_n_49_0));
  INV_X1_LVT execution_unit_0_i_44_0 (.ZN(execution_unit_0_n_44_0), .A(
      e_state[2]));
  NAND4_X1_LVT execution_unit_0_i_44_1 (.ZN(execution_unit_0_n_44_1), .A1(
      execution_unit_0_n_44_0), .A2(e_state[0]), .A3(e_state[1]), .A4(e_state[3]));
  DFFR_X1_LVT execution_unit_0_mdb_in_buf_en_reg (.Q(
      execution_unit_0_mdb_in_buf_en), .QN(), .CK(cpu_mclk), .D(
      execution_unit_0_n_1), .RN(execution_unit_0_n_18));
  AND2_X1_LVT execution_unit_0_i_44_2 (.ZN(execution_unit_0_n_96), .A1(
      execution_unit_0_n_44_1), .A2(execution_unit_0_mdb_in_buf_en));
  INV_X1_LVT execution_unit_0_i_45_0 (.ZN(execution_unit_0_n_45_0), .A(
      e_state[2]));
  NAND4_X1_LVT execution_unit_0_i_45_1 (.ZN(execution_unit_0_n_45_1), .A1(
      execution_unit_0_n_45_0), .A2(e_state[0]), .A3(e_state[1]), .A4(e_state[3]));
  NAND2_X1_LVT execution_unit_0_i_45_2 (.ZN(execution_unit_0_n_45_2), .A1(
      execution_unit_0_n_45_1), .A2(execution_unit_0_mdb_in_buf_en));
  NAND2_X1_LVT execution_unit_0_i_45_3 (.ZN(execution_unit_0_n_97), .A1(
      execution_unit_0_n_45_2), .A2(execution_unit_0_n_45_1));
  CLKGATETST_X1_LVT execution_unit_0_clk_gate_mdb_in_buf_valid_reg (.GCK(
      execution_unit_0_n_95), .CK(cpu_mclk), .E(execution_unit_0_n_97), .SE(1'b0));
  DFFR_X1_LVT execution_unit_0_mdb_in_buf_valid_reg (.Q(
      execution_unit_0_mdb_in_buf_valid), .QN(), .CK(execution_unit_0_n_95), .D(
      execution_unit_0_n_96), .RN(execution_unit_0_n_18));
  OAI21_X1_LVT execution_unit_0_i_48_5 (.ZN(execution_unit_0_n_48_3), .A(
      execution_unit_0_n_0), .B1(execution_unit_0_n_41), .B2(
      execution_unit_0_n_69));
  AND2_X1_LVT execution_unit_0_i_31_0 (.ZN(execution_unit_0_reg_sr_wr), .A1(
      execution_unit_0_n_4), .A2(inst_so[6]));
  INV_X1_LVT execution_unit_0_i_48_6 (.ZN(execution_unit_0_n_48_4), .A(
      execution_unit_0_reg_sr_wr));
  NAND2_X1_LVT execution_unit_0_i_48_7 (.ZN(execution_unit_0_n_101), .A1(
      execution_unit_0_n_48_3), .A2(execution_unit_0_n_48_4));
  NAND2_X1_LVT execution_unit_0_i_49_1 (.ZN(execution_unit_0_n_49_1), .A1(
      execution_unit_0_mdb_in_buf_valid), .A2(execution_unit_0_n_101));
  NOR2_X1_LVT execution_unit_0_i_49_9 (.ZN(execution_unit_0_n_105), .A1(
      execution_unit_0_n_49_7), .A2(execution_unit_0_n_49_1));
  CLKGATETST_X1_LVT execution_unit_0_clk_gate_mdb_in_buf_reg (.GCK(
      execution_unit_0_n_94), .CK(cpu_mclk), .E(execution_unit_0_mdb_in_buf_en), 
      .SE(1'b0));
  DFFR_X1_LVT \execution_unit_0_mdb_in_buf_reg[15] (.Q(
      execution_unit_0_mdb_in_buf[15]), .QN(), .CK(execution_unit_0_n_94), .D(
      execution_unit_0_n_65), .RN(execution_unit_0_n_18));
  NAND2_X1_LVT execution_unit_0_i_50_105 (.ZN(execution_unit_0_n_50_90), .A1(
      execution_unit_0_n_105), .A2(execution_unit_0_mdb_in_buf[15]));
  NAND2_X1_LVT execution_unit_0_i_49_2 (.ZN(execution_unit_0_n_49_2), .A1(
      execution_unit_0_n_49_0), .A2(execution_unit_0_n_49_1));
  INV_X1_LVT execution_unit_0_i_49_10 (.ZN(execution_unit_0_n_49_8), .A(
      execution_unit_0_n_101));
  NOR2_X1_LVT execution_unit_0_i_49_11 (.ZN(execution_unit_0_n_106), .A1(
      execution_unit_0_n_49_2), .A2(execution_unit_0_n_49_8));
  NAND2_X1_LVT execution_unit_0_i_50_106 (.ZN(execution_unit_0_n_50_91), .A1(
      execution_unit_0_n_106), .A2(execution_unit_0_n_65));
  NOR2_X1_LVT execution_unit_0_i_49_3 (.ZN(execution_unit_0_n_49_3), .A1(
      execution_unit_0_n_49_2), .A2(execution_unit_0_n_101));
  INV_X1_LVT execution_unit_0_i_20_0 (.ZN(execution_unit_0_n_39), .A(
      execution_unit_0_n_38));
  NAND2_X1_LVT execution_unit_0_i_48_2 (.ZN(execution_unit_0_n_48_1), .A1(
      execution_unit_0_n_3), .A2(execution_unit_0_n_39));
  INV_X1_LVT execution_unit_0_i_48_3 (.ZN(execution_unit_0_n_48_2), .A(
      execution_unit_0_n_4));
  OAI21_X1_LVT execution_unit_0_i_48_4 (.ZN(execution_unit_0_n_100), .A(
      execution_unit_0_n_48_1), .B1(execution_unit_0_n_48_2), .B2(
      execution_unit_0_n_37));
  AND2_X1_LVT execution_unit_0_i_49_12 (.ZN(execution_unit_0_n_107), .A1(
      execution_unit_0_n_49_3), .A2(execution_unit_0_n_100));
  NAND2_X1_LVT execution_unit_0_i_50_107 (.ZN(execution_unit_0_n_50_92), .A1(
      execution_unit_0_n_107), .A2(inst_dext[15]));
  INV_X1_LVT execution_unit_0_i_49_4 (.ZN(execution_unit_0_n_49_4), .A(
      execution_unit_0_n_100));
  NAND2_X1_LVT execution_unit_0_i_49_5 (.ZN(execution_unit_0_n_49_5), .A1(
      execution_unit_0_n_49_3), .A2(execution_unit_0_n_49_4));
  OR4_X1_LVT execution_unit_0_i_48_0 (.ZN(execution_unit_0_n_48_0), .A1(
      inst_as[7]), .A2(inst_as[5]), .A3(inst_type[1]), .A4(inst_so[6]));
  AND2_X1_LVT execution_unit_0_i_48_1 (.ZN(execution_unit_0_n_99), .A1(
      execution_unit_0_n_48_0), .A2(execution_unit_0_n_0));
  INV_X1_LVT execution_unit_0_i_49_13 (.ZN(execution_unit_0_n_49_9), .A(
      execution_unit_0_n_99));
  NOR2_X1_LVT execution_unit_0_i_49_14 (.ZN(execution_unit_0_n_108), .A1(
      execution_unit_0_n_49_5), .A2(execution_unit_0_n_49_9));
  NAND2_X1_LVT execution_unit_0_i_50_108 (.ZN(execution_unit_0_n_50_93), .A1(
      execution_unit_0_n_108), .A2(inst_sext[15]));
  NAND4_X1_LVT execution_unit_0_i_50_109 (.ZN(execution_unit_0_n_50_94), .A1(
      execution_unit_0_n_50_90), .A2(execution_unit_0_n_50_91), .A3(
      execution_unit_0_n_50_92), .A4(execution_unit_0_n_50_93));
  INV_X1_LVT execution_unit_0_i_49_6 (.ZN(execution_unit_0_n_49_6), .A(
      execution_unit_0_n_102));
  NOR2_X1_LVT execution_unit_0_i_49_7 (.ZN(execution_unit_0_n_104), .A1(
      execution_unit_0_n_49_6), .A2(execution_unit_0_n_103));
  AOI221_X1_LVT execution_unit_0_i_50_110 (.ZN(execution_unit_0_n_50_95), .A(
      execution_unit_0_n_50_94), .B1(execution_unit_0_n_103), .B2(
      execution_unit_0_reg_src[15]), .C1(execution_unit_0_n_104), .C2(
      dbg_reg_din[15]));
  INV_X1_LVT execution_unit_0_i_50_111 (.ZN(execution_unit_0_n_124), .A(
      execution_unit_0_n_50_95));
  DFFR_X1_LVT \execution_unit_0_mdb_in_buf_reg[14] (.Q(
      execution_unit_0_mdb_in_buf[14]), .QN(), .CK(execution_unit_0_n_94), .D(
      execution_unit_0_n_64), .RN(execution_unit_0_n_18));
  NAND2_X1_LVT execution_unit_0_i_50_98 (.ZN(execution_unit_0_n_50_84), .A1(
      execution_unit_0_n_105), .A2(execution_unit_0_mdb_in_buf[14]));
  NAND2_X1_LVT execution_unit_0_i_50_99 (.ZN(execution_unit_0_n_50_85), .A1(
      execution_unit_0_n_106), .A2(execution_unit_0_n_64));
  NAND2_X1_LVT execution_unit_0_i_50_100 (.ZN(execution_unit_0_n_50_86), .A1(
      execution_unit_0_n_107), .A2(inst_dext[14]));
  NAND2_X1_LVT execution_unit_0_i_50_101 (.ZN(execution_unit_0_n_50_87), .A1(
      execution_unit_0_n_108), .A2(inst_sext[14]));
  NAND4_X1_LVT execution_unit_0_i_50_102 (.ZN(execution_unit_0_n_50_88), .A1(
      execution_unit_0_n_50_84), .A2(execution_unit_0_n_50_85), .A3(
      execution_unit_0_n_50_86), .A4(execution_unit_0_n_50_87));
  AOI221_X1_LVT execution_unit_0_i_50_103 (.ZN(execution_unit_0_n_50_89), .A(
      execution_unit_0_n_50_88), .B1(execution_unit_0_n_103), .B2(
      execution_unit_0_reg_src[14]), .C1(execution_unit_0_n_104), .C2(
      dbg_reg_din[14]));
  INV_X1_LVT execution_unit_0_i_50_104 (.ZN(execution_unit_0_n_123), .A(
      execution_unit_0_n_50_89));
  DFFR_X1_LVT \execution_unit_0_mdb_in_buf_reg[13] (.Q(
      execution_unit_0_mdb_in_buf[13]), .QN(), .CK(execution_unit_0_n_94), .D(
      execution_unit_0_n_63), .RN(execution_unit_0_n_18));
  NAND2_X1_LVT execution_unit_0_i_50_91 (.ZN(execution_unit_0_n_50_78), .A1(
      execution_unit_0_n_105), .A2(execution_unit_0_mdb_in_buf[13]));
  NAND2_X1_LVT execution_unit_0_i_50_92 (.ZN(execution_unit_0_n_50_79), .A1(
      execution_unit_0_n_106), .A2(execution_unit_0_n_63));
  NAND2_X1_LVT execution_unit_0_i_50_93 (.ZN(execution_unit_0_n_50_80), .A1(
      execution_unit_0_n_107), .A2(inst_dext[13]));
  NAND2_X1_LVT execution_unit_0_i_50_94 (.ZN(execution_unit_0_n_50_81), .A1(
      execution_unit_0_n_108), .A2(inst_sext[13]));
  NAND4_X1_LVT execution_unit_0_i_50_95 (.ZN(execution_unit_0_n_50_82), .A1(
      execution_unit_0_n_50_78), .A2(execution_unit_0_n_50_79), .A3(
      execution_unit_0_n_50_80), .A4(execution_unit_0_n_50_81));
  AOI221_X1_LVT execution_unit_0_i_50_96 (.ZN(execution_unit_0_n_50_83), .A(
      execution_unit_0_n_50_82), .B1(execution_unit_0_n_103), .B2(
      execution_unit_0_reg_src[13]), .C1(execution_unit_0_n_104), .C2(
      dbg_reg_din[13]));
  INV_X1_LVT execution_unit_0_i_50_97 (.ZN(execution_unit_0_n_122), .A(
      execution_unit_0_n_50_83));
  DFFR_X1_LVT \execution_unit_0_mdb_in_buf_reg[12] (.Q(
      execution_unit_0_mdb_in_buf[12]), .QN(), .CK(execution_unit_0_n_94), .D(
      execution_unit_0_n_62), .RN(execution_unit_0_n_18));
  NAND2_X1_LVT execution_unit_0_i_50_84 (.ZN(execution_unit_0_n_50_72), .A1(
      execution_unit_0_n_105), .A2(execution_unit_0_mdb_in_buf[12]));
  NAND2_X1_LVT execution_unit_0_i_50_85 (.ZN(execution_unit_0_n_50_73), .A1(
      execution_unit_0_n_106), .A2(execution_unit_0_n_62));
  NAND2_X1_LVT execution_unit_0_i_50_86 (.ZN(execution_unit_0_n_50_74), .A1(
      execution_unit_0_n_107), .A2(inst_dext[12]));
  NAND2_X1_LVT execution_unit_0_i_50_87 (.ZN(execution_unit_0_n_50_75), .A1(
      execution_unit_0_n_108), .A2(inst_sext[12]));
  NAND4_X1_LVT execution_unit_0_i_50_88 (.ZN(execution_unit_0_n_50_76), .A1(
      execution_unit_0_n_50_72), .A2(execution_unit_0_n_50_73), .A3(
      execution_unit_0_n_50_74), .A4(execution_unit_0_n_50_75));
  AOI221_X1_LVT execution_unit_0_i_50_89 (.ZN(execution_unit_0_n_50_77), .A(
      execution_unit_0_n_50_76), .B1(execution_unit_0_n_103), .B2(
      execution_unit_0_reg_src[12]), .C1(execution_unit_0_n_104), .C2(
      dbg_reg_din[12]));
  INV_X1_LVT execution_unit_0_i_50_90 (.ZN(execution_unit_0_n_121), .A(
      execution_unit_0_n_50_77));
  DFFR_X1_LVT \execution_unit_0_mdb_in_buf_reg[11] (.Q(
      execution_unit_0_mdb_in_buf[11]), .QN(), .CK(execution_unit_0_n_94), .D(
      execution_unit_0_n_61), .RN(execution_unit_0_n_18));
  NAND2_X1_LVT execution_unit_0_i_50_77 (.ZN(execution_unit_0_n_50_66), .A1(
      execution_unit_0_n_105), .A2(execution_unit_0_mdb_in_buf[11]));
  NAND2_X1_LVT execution_unit_0_i_50_78 (.ZN(execution_unit_0_n_50_67), .A1(
      execution_unit_0_n_106), .A2(execution_unit_0_n_61));
  NAND2_X1_LVT execution_unit_0_i_50_79 (.ZN(execution_unit_0_n_50_68), .A1(
      execution_unit_0_n_107), .A2(inst_dext[11]));
  NAND2_X1_LVT execution_unit_0_i_50_80 (.ZN(execution_unit_0_n_50_69), .A1(
      execution_unit_0_n_108), .A2(inst_sext[11]));
  NAND4_X1_LVT execution_unit_0_i_50_81 (.ZN(execution_unit_0_n_50_70), .A1(
      execution_unit_0_n_50_66), .A2(execution_unit_0_n_50_67), .A3(
      execution_unit_0_n_50_68), .A4(execution_unit_0_n_50_69));
  AOI221_X1_LVT execution_unit_0_i_50_82 (.ZN(execution_unit_0_n_50_71), .A(
      execution_unit_0_n_50_70), .B1(execution_unit_0_n_103), .B2(
      execution_unit_0_reg_src[11]), .C1(execution_unit_0_n_104), .C2(
      dbg_reg_din[11]));
  INV_X1_LVT execution_unit_0_i_50_83 (.ZN(execution_unit_0_n_120), .A(
      execution_unit_0_n_50_71));
  DFFR_X1_LVT \execution_unit_0_mdb_in_buf_reg[10] (.Q(
      execution_unit_0_mdb_in_buf[10]), .QN(), .CK(execution_unit_0_n_94), .D(
      execution_unit_0_n_60), .RN(execution_unit_0_n_18));
  NAND2_X1_LVT execution_unit_0_i_50_70 (.ZN(execution_unit_0_n_50_60), .A1(
      execution_unit_0_n_105), .A2(execution_unit_0_mdb_in_buf[10]));
  NAND2_X1_LVT execution_unit_0_i_50_71 (.ZN(execution_unit_0_n_50_61), .A1(
      execution_unit_0_n_106), .A2(execution_unit_0_n_60));
  NAND2_X1_LVT execution_unit_0_i_50_72 (.ZN(execution_unit_0_n_50_62), .A1(
      execution_unit_0_n_107), .A2(inst_dext[10]));
  NAND2_X1_LVT execution_unit_0_i_50_73 (.ZN(execution_unit_0_n_50_63), .A1(
      execution_unit_0_n_108), .A2(inst_sext[10]));
  NAND4_X1_LVT execution_unit_0_i_50_74 (.ZN(execution_unit_0_n_50_64), .A1(
      execution_unit_0_n_50_60), .A2(execution_unit_0_n_50_61), .A3(
      execution_unit_0_n_50_62), .A4(execution_unit_0_n_50_63));
  AOI221_X1_LVT execution_unit_0_i_50_75 (.ZN(execution_unit_0_n_50_65), .A(
      execution_unit_0_n_50_64), .B1(execution_unit_0_n_103), .B2(
      execution_unit_0_reg_src[10]), .C1(execution_unit_0_n_104), .C2(
      dbg_reg_din[10]));
  INV_X1_LVT execution_unit_0_i_50_76 (.ZN(execution_unit_0_n_119), .A(
      execution_unit_0_n_50_65));
  DFFR_X1_LVT \execution_unit_0_mdb_in_buf_reg[9] (.Q(
      execution_unit_0_mdb_in_buf[9]), .QN(), .CK(execution_unit_0_n_94), .D(
      execution_unit_0_n_59), .RN(execution_unit_0_n_18));
  NAND2_X1_LVT execution_unit_0_i_50_63 (.ZN(execution_unit_0_n_50_54), .A1(
      execution_unit_0_n_105), .A2(execution_unit_0_mdb_in_buf[9]));
  NAND2_X1_LVT execution_unit_0_i_50_64 (.ZN(execution_unit_0_n_50_55), .A1(
      execution_unit_0_n_106), .A2(execution_unit_0_n_59));
  NAND2_X1_LVT execution_unit_0_i_50_65 (.ZN(execution_unit_0_n_50_56), .A1(
      execution_unit_0_n_107), .A2(inst_dext[9]));
  NAND2_X1_LVT execution_unit_0_i_50_66 (.ZN(execution_unit_0_n_50_57), .A1(
      execution_unit_0_n_108), .A2(inst_sext[9]));
  NAND4_X1_LVT execution_unit_0_i_50_67 (.ZN(execution_unit_0_n_50_58), .A1(
      execution_unit_0_n_50_54), .A2(execution_unit_0_n_50_55), .A3(
      execution_unit_0_n_50_56), .A4(execution_unit_0_n_50_57));
  AOI221_X1_LVT execution_unit_0_i_50_68 (.ZN(execution_unit_0_n_50_59), .A(
      execution_unit_0_n_50_58), .B1(execution_unit_0_n_103), .B2(
      execution_unit_0_reg_src[9]), .C1(execution_unit_0_n_104), .C2(
      dbg_reg_din[9]));
  INV_X1_LVT execution_unit_0_i_50_69 (.ZN(execution_unit_0_n_118), .A(
      execution_unit_0_n_50_59));
  DFFR_X1_LVT \execution_unit_0_mdb_in_buf_reg[8] (.Q(
      execution_unit_0_mdb_in_buf[8]), .QN(), .CK(execution_unit_0_n_94), .D(
      execution_unit_0_n_58), .RN(execution_unit_0_n_18));
  NAND2_X1_LVT execution_unit_0_i_50_56 (.ZN(execution_unit_0_n_50_48), .A1(
      execution_unit_0_n_105), .A2(execution_unit_0_mdb_in_buf[8]));
  NAND2_X1_LVT execution_unit_0_i_50_57 (.ZN(execution_unit_0_n_50_49), .A1(
      execution_unit_0_n_106), .A2(execution_unit_0_n_58));
  NAND2_X1_LVT execution_unit_0_i_50_58 (.ZN(execution_unit_0_n_50_50), .A1(
      execution_unit_0_n_107), .A2(inst_dext[8]));
  NAND2_X1_LVT execution_unit_0_i_50_59 (.ZN(execution_unit_0_n_50_51), .A1(
      execution_unit_0_n_108), .A2(inst_sext[8]));
  NAND4_X1_LVT execution_unit_0_i_50_60 (.ZN(execution_unit_0_n_50_52), .A1(
      execution_unit_0_n_50_48), .A2(execution_unit_0_n_50_49), .A3(
      execution_unit_0_n_50_50), .A4(execution_unit_0_n_50_51));
  AOI221_X1_LVT execution_unit_0_i_50_61 (.ZN(execution_unit_0_n_50_53), .A(
      execution_unit_0_n_50_52), .B1(execution_unit_0_n_103), .B2(
      execution_unit_0_reg_src[8]), .C1(execution_unit_0_n_104), .C2(
      dbg_reg_din[8]));
  INV_X1_LVT execution_unit_0_i_50_62 (.ZN(execution_unit_0_n_117), .A(
      execution_unit_0_n_50_53));
  DFFR_X1_LVT \execution_unit_0_mdb_in_buf_reg[7] (.Q(
      execution_unit_0_mdb_in_buf[7]), .QN(), .CK(execution_unit_0_n_94), .D(
      execution_unit_0_n_57), .RN(execution_unit_0_n_18));
  NAND2_X1_LVT execution_unit_0_i_50_49 (.ZN(execution_unit_0_n_50_42), .A1(
      execution_unit_0_n_105), .A2(execution_unit_0_mdb_in_buf[7]));
  NAND2_X1_LVT execution_unit_0_i_50_50 (.ZN(execution_unit_0_n_50_43), .A1(
      execution_unit_0_n_106), .A2(execution_unit_0_n_57));
  NAND2_X1_LVT execution_unit_0_i_50_51 (.ZN(execution_unit_0_n_50_44), .A1(
      execution_unit_0_n_107), .A2(inst_dext[7]));
  NAND2_X1_LVT execution_unit_0_i_50_52 (.ZN(execution_unit_0_n_50_45), .A1(
      execution_unit_0_n_108), .A2(inst_sext[7]));
  NAND4_X1_LVT execution_unit_0_i_50_53 (.ZN(execution_unit_0_n_50_46), .A1(
      execution_unit_0_n_50_42), .A2(execution_unit_0_n_50_43), .A3(
      execution_unit_0_n_50_44), .A4(execution_unit_0_n_50_45));
  AOI221_X1_LVT execution_unit_0_i_50_54 (.ZN(execution_unit_0_n_50_47), .A(
      execution_unit_0_n_50_46), .B1(execution_unit_0_n_103), .B2(
      execution_unit_0_reg_src[7]), .C1(execution_unit_0_n_104), .C2(
      dbg_reg_din[7]));
  INV_X1_LVT execution_unit_0_i_50_55 (.ZN(execution_unit_0_n_116), .A(
      execution_unit_0_n_50_47));
  DFFR_X1_LVT \execution_unit_0_mdb_in_buf_reg[6] (.Q(
      execution_unit_0_mdb_in_buf[6]), .QN(), .CK(execution_unit_0_n_94), .D(
      execution_unit_0_n_56), .RN(execution_unit_0_n_18));
  NAND2_X1_LVT execution_unit_0_i_50_42 (.ZN(execution_unit_0_n_50_36), .A1(
      execution_unit_0_n_105), .A2(execution_unit_0_mdb_in_buf[6]));
  NAND2_X1_LVT execution_unit_0_i_50_43 (.ZN(execution_unit_0_n_50_37), .A1(
      execution_unit_0_n_106), .A2(execution_unit_0_n_56));
  NAND2_X1_LVT execution_unit_0_i_50_44 (.ZN(execution_unit_0_n_50_38), .A1(
      execution_unit_0_n_107), .A2(inst_dext[6]));
  NAND2_X1_LVT execution_unit_0_i_50_45 (.ZN(execution_unit_0_n_50_39), .A1(
      execution_unit_0_n_108), .A2(inst_sext[6]));
  NAND4_X1_LVT execution_unit_0_i_50_46 (.ZN(execution_unit_0_n_50_40), .A1(
      execution_unit_0_n_50_36), .A2(execution_unit_0_n_50_37), .A3(
      execution_unit_0_n_50_38), .A4(execution_unit_0_n_50_39));
  AOI221_X1_LVT execution_unit_0_i_50_47 (.ZN(execution_unit_0_n_50_41), .A(
      execution_unit_0_n_50_40), .B1(execution_unit_0_n_103), .B2(
      execution_unit_0_reg_src[6]), .C1(execution_unit_0_n_104), .C2(
      dbg_reg_din[6]));
  INV_X1_LVT execution_unit_0_i_50_48 (.ZN(execution_unit_0_n_115), .A(
      execution_unit_0_n_50_41));
  DFFR_X1_LVT \execution_unit_0_mdb_in_buf_reg[5] (.Q(
      execution_unit_0_mdb_in_buf[5]), .QN(), .CK(execution_unit_0_n_94), .D(
      execution_unit_0_n_55), .RN(execution_unit_0_n_18));
  NAND2_X1_LVT execution_unit_0_i_50_35 (.ZN(execution_unit_0_n_50_30), .A1(
      execution_unit_0_n_105), .A2(execution_unit_0_mdb_in_buf[5]));
  NAND2_X1_LVT execution_unit_0_i_50_36 (.ZN(execution_unit_0_n_50_31), .A1(
      execution_unit_0_n_106), .A2(execution_unit_0_n_55));
  NAND2_X1_LVT execution_unit_0_i_50_37 (.ZN(execution_unit_0_n_50_32), .A1(
      execution_unit_0_n_107), .A2(inst_dext[5]));
  NAND2_X1_LVT execution_unit_0_i_50_38 (.ZN(execution_unit_0_n_50_33), .A1(
      execution_unit_0_n_108), .A2(inst_sext[5]));
  NAND4_X1_LVT execution_unit_0_i_50_39 (.ZN(execution_unit_0_n_50_34), .A1(
      execution_unit_0_n_50_30), .A2(execution_unit_0_n_50_31), .A3(
      execution_unit_0_n_50_32), .A4(execution_unit_0_n_50_33));
  AOI221_X1_LVT execution_unit_0_i_50_40 (.ZN(execution_unit_0_n_50_35), .A(
      execution_unit_0_n_50_34), .B1(execution_unit_0_n_103), .B2(
      execution_unit_0_reg_src[5]), .C1(execution_unit_0_n_104), .C2(
      dbg_reg_din[5]));
  INV_X1_LVT execution_unit_0_i_50_41 (.ZN(execution_unit_0_n_114), .A(
      execution_unit_0_n_50_35));
  DFFR_X1_LVT \execution_unit_0_mdb_in_buf_reg[4] (.Q(
      execution_unit_0_mdb_in_buf[4]), .QN(), .CK(execution_unit_0_n_94), .D(
      execution_unit_0_n_54), .RN(execution_unit_0_n_18));
  NAND2_X1_LVT execution_unit_0_i_50_28 (.ZN(execution_unit_0_n_50_24), .A1(
      execution_unit_0_n_105), .A2(execution_unit_0_mdb_in_buf[4]));
  NAND2_X1_LVT execution_unit_0_i_50_29 (.ZN(execution_unit_0_n_50_25), .A1(
      execution_unit_0_n_106), .A2(execution_unit_0_n_54));
  NAND2_X1_LVT execution_unit_0_i_50_30 (.ZN(execution_unit_0_n_50_26), .A1(
      execution_unit_0_n_107), .A2(inst_dext[4]));
  NAND2_X1_LVT execution_unit_0_i_50_31 (.ZN(execution_unit_0_n_50_27), .A1(
      execution_unit_0_n_108), .A2(inst_sext[4]));
  NAND4_X1_LVT execution_unit_0_i_50_32 (.ZN(execution_unit_0_n_50_28), .A1(
      execution_unit_0_n_50_24), .A2(execution_unit_0_n_50_25), .A3(
      execution_unit_0_n_50_26), .A4(execution_unit_0_n_50_27));
  AOI221_X1_LVT execution_unit_0_i_50_33 (.ZN(execution_unit_0_n_50_29), .A(
      execution_unit_0_n_50_28), .B1(execution_unit_0_n_103), .B2(
      execution_unit_0_reg_src[4]), .C1(execution_unit_0_n_104), .C2(
      dbg_reg_din[4]));
  INV_X1_LVT execution_unit_0_i_50_34 (.ZN(execution_unit_0_n_113), .A(
      execution_unit_0_n_50_29));
  DFFR_X1_LVT \execution_unit_0_mdb_in_buf_reg[3] (.Q(
      execution_unit_0_mdb_in_buf[3]), .QN(), .CK(execution_unit_0_n_94), .D(
      execution_unit_0_n_53), .RN(execution_unit_0_n_18));
  NAND2_X1_LVT execution_unit_0_i_50_21 (.ZN(execution_unit_0_n_50_18), .A1(
      execution_unit_0_n_105), .A2(execution_unit_0_mdb_in_buf[3]));
  NAND2_X1_LVT execution_unit_0_i_50_22 (.ZN(execution_unit_0_n_50_19), .A1(
      execution_unit_0_n_106), .A2(execution_unit_0_n_53));
  NAND2_X1_LVT execution_unit_0_i_50_23 (.ZN(execution_unit_0_n_50_20), .A1(
      execution_unit_0_n_107), .A2(inst_dext[3]));
  NAND2_X1_LVT execution_unit_0_i_50_24 (.ZN(execution_unit_0_n_50_21), .A1(
      execution_unit_0_n_108), .A2(inst_sext[3]));
  NAND4_X1_LVT execution_unit_0_i_50_25 (.ZN(execution_unit_0_n_50_22), .A1(
      execution_unit_0_n_50_18), .A2(execution_unit_0_n_50_19), .A3(
      execution_unit_0_n_50_20), .A4(execution_unit_0_n_50_21));
  AOI221_X1_LVT execution_unit_0_i_50_26 (.ZN(execution_unit_0_n_50_23), .A(
      execution_unit_0_n_50_22), .B1(execution_unit_0_n_103), .B2(
      execution_unit_0_reg_src[3]), .C1(execution_unit_0_n_104), .C2(
      dbg_reg_din[3]));
  INV_X1_LVT execution_unit_0_i_50_27 (.ZN(execution_unit_0_n_112), .A(
      execution_unit_0_n_50_23));
  DFFR_X1_LVT \execution_unit_0_mdb_in_buf_reg[2] (.Q(
      execution_unit_0_mdb_in_buf[2]), .QN(), .CK(execution_unit_0_n_94), .D(
      execution_unit_0_n_52), .RN(execution_unit_0_n_18));
  NAND2_X1_LVT execution_unit_0_i_50_14 (.ZN(execution_unit_0_n_50_12), .A1(
      execution_unit_0_n_105), .A2(execution_unit_0_mdb_in_buf[2]));
  NAND2_X1_LVT execution_unit_0_i_50_15 (.ZN(execution_unit_0_n_50_13), .A1(
      execution_unit_0_n_106), .A2(execution_unit_0_n_52));
  NAND2_X1_LVT execution_unit_0_i_50_16 (.ZN(execution_unit_0_n_50_14), .A1(
      execution_unit_0_n_107), .A2(inst_dext[2]));
  NAND2_X1_LVT execution_unit_0_i_50_17 (.ZN(execution_unit_0_n_50_15), .A1(
      execution_unit_0_n_108), .A2(inst_sext[2]));
  NAND4_X1_LVT execution_unit_0_i_50_18 (.ZN(execution_unit_0_n_50_16), .A1(
      execution_unit_0_n_50_12), .A2(execution_unit_0_n_50_13), .A3(
      execution_unit_0_n_50_14), .A4(execution_unit_0_n_50_15));
  AOI221_X1_LVT execution_unit_0_i_50_19 (.ZN(execution_unit_0_n_50_17), .A(
      execution_unit_0_n_50_16), .B1(execution_unit_0_n_103), .B2(
      execution_unit_0_reg_src[2]), .C1(execution_unit_0_n_104), .C2(
      dbg_reg_din[2]));
  INV_X1_LVT execution_unit_0_i_50_20 (.ZN(execution_unit_0_n_111), .A(
      execution_unit_0_n_50_17));
  DFFR_X1_LVT \execution_unit_0_mdb_in_buf_reg[1] (.Q(
      execution_unit_0_mdb_in_buf[1]), .QN(), .CK(execution_unit_0_n_94), .D(
      execution_unit_0_n_51), .RN(execution_unit_0_n_18));
  NAND2_X1_LVT execution_unit_0_i_50_7 (.ZN(execution_unit_0_n_50_6), .A1(
      execution_unit_0_n_105), .A2(execution_unit_0_mdb_in_buf[1]));
  NAND2_X1_LVT execution_unit_0_i_50_8 (.ZN(execution_unit_0_n_50_7), .A1(
      execution_unit_0_n_106), .A2(execution_unit_0_n_51));
  NAND2_X1_LVT execution_unit_0_i_50_9 (.ZN(execution_unit_0_n_50_8), .A1(
      execution_unit_0_n_107), .A2(inst_dext[1]));
  NAND2_X1_LVT execution_unit_0_i_50_10 (.ZN(execution_unit_0_n_50_9), .A1(
      execution_unit_0_n_108), .A2(inst_sext[1]));
  NAND4_X1_LVT execution_unit_0_i_50_11 (.ZN(execution_unit_0_n_50_10), .A1(
      execution_unit_0_n_50_6), .A2(execution_unit_0_n_50_7), .A3(
      execution_unit_0_n_50_8), .A4(execution_unit_0_n_50_9));
  AOI221_X1_LVT execution_unit_0_i_50_12 (.ZN(execution_unit_0_n_50_11), .A(
      execution_unit_0_n_50_10), .B1(execution_unit_0_n_103), .B2(
      execution_unit_0_reg_src[1]), .C1(execution_unit_0_n_104), .C2(
      dbg_reg_din[1]));
  INV_X1_LVT execution_unit_0_i_50_13 (.ZN(execution_unit_0_n_110), .A(
      execution_unit_0_n_50_11));
  DFFR_X1_LVT \execution_unit_0_mdb_in_buf_reg[0] (.Q(
      execution_unit_0_mdb_in_buf[0]), .QN(), .CK(execution_unit_0_n_94), .D(
      execution_unit_0_n_50), .RN(execution_unit_0_n_18));
  NAND2_X1_LVT execution_unit_0_i_50_0 (.ZN(execution_unit_0_n_50_0), .A1(
      execution_unit_0_mdb_in_buf[0]), .A2(execution_unit_0_n_105));
  NAND2_X1_LVT execution_unit_0_i_50_1 (.ZN(execution_unit_0_n_50_1), .A1(
      execution_unit_0_n_50), .A2(execution_unit_0_n_106));
  NAND2_X1_LVT execution_unit_0_i_50_2 (.ZN(execution_unit_0_n_50_2), .A1(
      inst_dext[0]), .A2(execution_unit_0_n_107));
  NAND2_X1_LVT execution_unit_0_i_50_3 (.ZN(execution_unit_0_n_50_3), .A1(
      inst_sext[0]), .A2(execution_unit_0_n_108));
  NAND4_X1_LVT execution_unit_0_i_50_4 (.ZN(execution_unit_0_n_50_4), .A1(
      execution_unit_0_n_50_0), .A2(execution_unit_0_n_50_1), .A3(
      execution_unit_0_n_50_2), .A4(execution_unit_0_n_50_3));
  AOI221_X1_LVT execution_unit_0_i_50_5 (.ZN(execution_unit_0_n_50_5), .A(
      execution_unit_0_n_50_4), .B1(execution_unit_0_reg_src[0]), .B2(
      execution_unit_0_n_103), .C1(dbg_reg_din[0]), .C2(execution_unit_0_n_104));
  INV_X1_LVT execution_unit_0_i_50_6 (.ZN(execution_unit_0_n_109), .A(
      execution_unit_0_n_50_5));
  OR3_X1_LVT execution_unit_0_alu_0_i_42_0 (.ZN(execution_unit_0_alu_0_n_104), 
      .A1(inst_so[7]), .A2(inst_alu[3]), .A3(cpu_halt_st));
  NAND2_X1_LVT execution_unit_0_alu_0_i_0_0 (.ZN(
      execution_unit_0_alu_0_op_bit8_msk), .A1(execution_unit_0_n_0), .A2(
      inst_bw));
  AND2_X1_LVT execution_unit_0_alu_0_i_1_7 (.ZN(execution_unit_0_alu_0_n_7), .A1(
      execution_unit_0_alu_0_op_bit8_msk), .A2(execution_unit_0_n_93));
  XOR2_X1_LVT execution_unit_0_alu_0_i_29_0 (.Z(execution_unit_0_alu_0_n_86), .A(
      execution_unit_0_status[3]), .B(execution_unit_0_status[2]));
  INV_X1_LVT execution_unit_0_alu_0_i_30_0 (.ZN(execution_unit_0_alu_0_n_30_0), 
      .A(execution_unit_0_alu_0_n_86));
  INV_X1_LVT execution_unit_0_alu_0_i_30_1 (.ZN(execution_unit_0_alu_0_n_30_1), 
      .A(execution_unit_0_status[1]));
  INV_X1_LVT execution_unit_0_alu_0_i_30_2 (.ZN(execution_unit_0_alu_0_n_30_2), 
      .A(execution_unit_0_status[0]));
  AOI222_X1_LVT execution_unit_0_alu_0_i_30_3 (.ZN(execution_unit_0_alu_0_n_30_3), 
      .A1(execution_unit_0_alu_0_n_30_0), .A2(inst_jmp[6]), .B1(
      execution_unit_0_alu_0_n_30_1), .B2(inst_jmp[1]), .C1(
      execution_unit_0_alu_0_n_30_2), .C2(inst_jmp[3]));
  INV_X1_LVT execution_unit_0_alu_0_i_30_4 (.ZN(execution_unit_0_alu_0_n_30_4), 
      .A(execution_unit_0_status[2]));
  NAND2_X1_LVT execution_unit_0_alu_0_i_30_5 (.ZN(execution_unit_0_alu_0_n_30_5), 
      .A1(execution_unit_0_alu_0_n_30_4), .A2(inst_jmp[4]));
  NAND2_X1_LVT execution_unit_0_alu_0_i_30_6 (.ZN(execution_unit_0_alu_0_n_30_6), 
      .A1(inst_jmp[0]), .A2(execution_unit_0_status[1]));
  NAND2_X1_LVT execution_unit_0_alu_0_i_30_7 (.ZN(execution_unit_0_alu_0_n_30_7), 
      .A1(inst_jmp[2]), .A2(execution_unit_0_status[0]));
  NAND2_X1_LVT execution_unit_0_alu_0_i_30_8 (.ZN(execution_unit_0_alu_0_n_30_8), 
      .A1(execution_unit_0_alu_0_n_86), .A2(inst_jmp[5]));
  AND4_X1_LVT execution_unit_0_alu_0_i_30_9 (.ZN(execution_unit_0_alu_0_n_30_9), 
      .A1(execution_unit_0_alu_0_n_30_5), .A2(execution_unit_0_alu_0_n_30_6), 
      .A3(execution_unit_0_alu_0_n_30_7), .A4(execution_unit_0_alu_0_n_30_8));
  AND2_X1_LVT execution_unit_0_alu_0_i_30_10 (.ZN(execution_unit_0_alu_0_n_87), 
      .A1(execution_unit_0_alu_0_n_30_3), .A2(execution_unit_0_alu_0_n_30_9));
  AND2_X1_LVT execution_unit_0_alu_0_i_2_0 (.ZN(
      execution_unit_0_alu_0_op_src_inv_cmd), .A1(execution_unit_0_n_0), .A2(
      inst_alu[0]));
  XNOR2_X1_LVT execution_unit_0_alu_0_i_4_15 (.ZN(execution_unit_0_alu_0_n_4_8), 
      .A(execution_unit_0_alu_0_op_src_inv_cmd), .B(execution_unit_0_n_124));
  INV_X1_LVT execution_unit_0_alu_0_i_4_1 (.ZN(execution_unit_0_alu_0_n_4_1), .A(
      execution_unit_0_alu_0_op_bit8_msk));
  NOR2_X1_LVT execution_unit_0_alu_0_i_4_16 (.ZN(execution_unit_0_alu_0_X[3]), 
      .A1(execution_unit_0_alu_0_n_4_8), .A2(execution_unit_0_alu_0_n_4_1));
  AND2_X1_LVT execution_unit_0_alu_0_i_39_7 (.ZN(execution_unit_0_alu_0_n_103), 
      .A1(execution_unit_0_alu_0_n_87), .A2(execution_unit_0_alu_0_X[3]));
  AND2_X1_LVT execution_unit_0_alu_0_i_1_6 (.ZN(execution_unit_0_alu_0_n_6), .A1(
      execution_unit_0_alu_0_op_bit8_msk), .A2(execution_unit_0_n_92));
  XNOR2_X1_LVT execution_unit_0_alu_0_i_4_13 (.ZN(execution_unit_0_alu_0_n_4_7), 
      .A(execution_unit_0_alu_0_op_src_inv_cmd), .B(execution_unit_0_n_123));
  NOR2_X1_LVT execution_unit_0_alu_0_i_4_14 (.ZN(execution_unit_0_alu_0_X[2]), 
      .A1(execution_unit_0_alu_0_n_4_7), .A2(execution_unit_0_alu_0_n_4_1));
  AND2_X1_LVT execution_unit_0_alu_0_i_39_6 (.ZN(execution_unit_0_alu_0_n_102), 
      .A1(execution_unit_0_alu_0_n_87), .A2(execution_unit_0_alu_0_X[2]));
  AND2_X1_LVT execution_unit_0_alu_0_i_1_5 (.ZN(execution_unit_0_alu_0_n_5), .A1(
      execution_unit_0_alu_0_op_bit8_msk), .A2(execution_unit_0_n_91));
  XNOR2_X1_LVT execution_unit_0_alu_0_i_4_11 (.ZN(execution_unit_0_alu_0_n_4_6), 
      .A(execution_unit_0_alu_0_op_src_inv_cmd), .B(execution_unit_0_n_122));
  NOR2_X1_LVT execution_unit_0_alu_0_i_4_12 (.ZN(execution_unit_0_alu_0_X[1]), 
      .A1(execution_unit_0_alu_0_n_4_6), .A2(execution_unit_0_alu_0_n_4_1));
  AND2_X1_LVT execution_unit_0_alu_0_i_39_5 (.ZN(execution_unit_0_alu_0_n_101), 
      .A1(execution_unit_0_alu_0_n_87), .A2(execution_unit_0_alu_0_X[1]));
  AND2_X1_LVT execution_unit_0_alu_0_i_1_4 (.ZN(execution_unit_0_alu_0_n_4), .A1(
      execution_unit_0_alu_0_op_bit8_msk), .A2(execution_unit_0_n_90));
  XNOR2_X1_LVT execution_unit_0_alu_0_i_4_9 (.ZN(execution_unit_0_alu_0_n_4_5), 
      .A(execution_unit_0_alu_0_op_src_inv_cmd), .B(execution_unit_0_n_121));
  NOR2_X1_LVT execution_unit_0_alu_0_i_4_10 (.ZN(execution_unit_0_alu_0_X[0]), 
      .A1(execution_unit_0_alu_0_n_4_5), .A2(execution_unit_0_alu_0_n_4_1));
  AND2_X1_LVT execution_unit_0_alu_0_i_39_4 (.ZN(execution_unit_0_alu_0_n_100), 
      .A1(execution_unit_0_alu_0_n_87), .A2(execution_unit_0_alu_0_X[0]));
  AND2_X1_LVT execution_unit_0_alu_0_i_1_3 (.ZN(execution_unit_0_alu_0_n_3), .A1(
      execution_unit_0_alu_0_op_bit8_msk), .A2(execution_unit_0_n_89));
  XNOR2_X1_LVT execution_unit_0_alu_0_i_4_7 (.ZN(execution_unit_0_alu_0_n_4_4), 
      .A(execution_unit_0_alu_0_op_src_inv_cmd), .B(execution_unit_0_n_120));
  NOR2_X1_LVT execution_unit_0_alu_0_i_4_8 (.ZN(execution_unit_0_alu_0_n_19), 
      .A1(execution_unit_0_alu_0_n_4_4), .A2(execution_unit_0_alu_0_n_4_1));
  AND2_X1_LVT execution_unit_0_alu_0_i_39_3 (.ZN(execution_unit_0_alu_0_n_99), 
      .A1(execution_unit_0_alu_0_n_87), .A2(execution_unit_0_alu_0_n_19));
  AND2_X1_LVT execution_unit_0_alu_0_i_1_2 (.ZN(execution_unit_0_alu_0_n_2), .A1(
      execution_unit_0_alu_0_op_bit8_msk), .A2(execution_unit_0_n_88));
  XNOR2_X1_LVT execution_unit_0_alu_0_i_4_5 (.ZN(execution_unit_0_alu_0_n_4_3), 
      .A(execution_unit_0_alu_0_op_src_inv_cmd), .B(execution_unit_0_n_119));
  NOR2_X1_LVT execution_unit_0_alu_0_i_4_6 (.ZN(execution_unit_0_alu_0_n_18), 
      .A1(execution_unit_0_alu_0_n_4_3), .A2(execution_unit_0_alu_0_n_4_1));
  AND2_X1_LVT execution_unit_0_alu_0_i_39_2 (.ZN(execution_unit_0_alu_0_n_98), 
      .A1(execution_unit_0_alu_0_n_87), .A2(execution_unit_0_alu_0_n_18));
  AND2_X1_LVT execution_unit_0_alu_0_i_1_1 (.ZN(execution_unit_0_alu_0_n_1), .A1(
      execution_unit_0_alu_0_op_bit8_msk), .A2(execution_unit_0_n_87));
  XNOR2_X1_LVT execution_unit_0_alu_0_i_4_3 (.ZN(execution_unit_0_alu_0_n_4_2), 
      .A(execution_unit_0_alu_0_op_src_inv_cmd), .B(execution_unit_0_n_118));
  NOR2_X1_LVT execution_unit_0_alu_0_i_4_4 (.ZN(execution_unit_0_alu_0_n_17), 
      .A1(execution_unit_0_alu_0_n_4_2), .A2(execution_unit_0_alu_0_n_4_1));
  AND2_X1_LVT execution_unit_0_alu_0_i_39_1 (.ZN(execution_unit_0_alu_0_n_97), 
      .A1(execution_unit_0_alu_0_n_87), .A2(execution_unit_0_alu_0_n_17));
  AND2_X1_LVT execution_unit_0_alu_0_i_1_0 (.ZN(execution_unit_0_alu_0_n_0), .A1(
      execution_unit_0_n_86), .A2(execution_unit_0_alu_0_op_bit8_msk));
  XNOR2_X1_LVT execution_unit_0_alu_0_i_4_0 (.ZN(execution_unit_0_alu_0_n_4_0), 
      .A(execution_unit_0_alu_0_op_src_inv_cmd), .B(execution_unit_0_n_117));
  NOR2_X1_LVT execution_unit_0_alu_0_i_4_2 (.ZN(execution_unit_0_alu_0_n_16), 
      .A1(execution_unit_0_alu_0_n_4_0), .A2(execution_unit_0_alu_0_n_4_1));
  AND2_X1_LVT execution_unit_0_alu_0_i_39_0 (.ZN(execution_unit_0_alu_0_n_96), 
      .A1(execution_unit_0_alu_0_n_16), .A2(execution_unit_0_alu_0_n_87));
  XOR2_X1_LVT execution_unit_0_alu_0_i_3_7 (.Z(execution_unit_0_alu_0_n_15), .A(
      execution_unit_0_alu_0_op_src_inv_cmd), .B(execution_unit_0_n_116));
  AND2_X1_LVT execution_unit_0_alu_0_i_38_0 (.ZN(execution_unit_0_alu_0_n_95), 
      .A1(execution_unit_0_alu_0_n_15), .A2(execution_unit_0_alu_0_n_87));
  XOR2_X1_LVT execution_unit_0_alu_0_i_3_6 (.Z(execution_unit_0_alu_0_n_14), .A(
      execution_unit_0_alu_0_op_src_inv_cmd), .B(execution_unit_0_n_115));
  AND2_X1_LVT execution_unit_0_alu_0_i_37_0 (.ZN(execution_unit_0_alu_0_n_94), 
      .A1(execution_unit_0_alu_0_n_14), .A2(execution_unit_0_alu_0_n_87));
  XOR2_X1_LVT execution_unit_0_alu_0_i_3_5 (.Z(execution_unit_0_alu_0_n_13), .A(
      execution_unit_0_alu_0_op_src_inv_cmd), .B(execution_unit_0_n_114));
  AND2_X1_LVT execution_unit_0_alu_0_i_36_0 (.ZN(execution_unit_0_alu_0_n_93), 
      .A1(execution_unit_0_alu_0_n_13), .A2(execution_unit_0_alu_0_n_87));
  XOR2_X1_LVT execution_unit_0_alu_0_i_3_4 (.Z(execution_unit_0_alu_0_n_12), .A(
      execution_unit_0_alu_0_op_src_inv_cmd), .B(execution_unit_0_n_113));
  AND2_X1_LVT execution_unit_0_alu_0_i_35_0 (.ZN(execution_unit_0_alu_0_n_92), 
      .A1(execution_unit_0_alu_0_n_12), .A2(execution_unit_0_alu_0_n_87));
  XOR2_X1_LVT execution_unit_0_alu_0_i_3_3 (.Z(execution_unit_0_alu_0_n_11), .A(
      execution_unit_0_alu_0_op_src_inv_cmd), .B(execution_unit_0_n_112));
  AND2_X1_LVT execution_unit_0_alu_0_i_34_0 (.ZN(execution_unit_0_alu_0_n_91), 
      .A1(execution_unit_0_alu_0_n_11), .A2(execution_unit_0_alu_0_n_87));
  XOR2_X1_LVT execution_unit_0_alu_0_i_3_2 (.Z(execution_unit_0_alu_0_n_10), .A(
      execution_unit_0_alu_0_op_src_inv_cmd), .B(execution_unit_0_n_111));
  AND2_X1_LVT execution_unit_0_alu_0_i_33_0 (.ZN(execution_unit_0_alu_0_n_90), 
      .A1(execution_unit_0_alu_0_n_10), .A2(execution_unit_0_alu_0_n_87));
  XOR2_X1_LVT execution_unit_0_alu_0_i_3_1 (.Z(execution_unit_0_alu_0_n_9), .A(
      execution_unit_0_alu_0_op_src_inv_cmd), .B(execution_unit_0_n_110));
  AND2_X1_LVT execution_unit_0_alu_0_i_32_0 (.ZN(execution_unit_0_alu_0_n_89), 
      .A1(execution_unit_0_alu_0_n_9), .A2(execution_unit_0_alu_0_n_87));
  XOR2_X1_LVT execution_unit_0_alu_0_i_3_0 (.Z(execution_unit_0_alu_0_n_8), .A(
      execution_unit_0_alu_0_op_src_inv_cmd), .B(execution_unit_0_n_109));
  AND2_X1_LVT execution_unit_0_alu_0_i_31_0 (.ZN(execution_unit_0_alu_0_n_88), 
      .A1(execution_unit_0_alu_0_n_8), .A2(execution_unit_0_alu_0_n_87));
  HA_X1_LVT execution_unit_0_alu_0_i_40_0 (.CO(execution_unit_0_alu_0_n_40_0), 
      .S(eu_mab[0]), .A(execution_unit_0_n_78), .B(execution_unit_0_alu_0_n_88));
  FA_X1_LVT execution_unit_0_alu_0_i_40_1 (.CO(execution_unit_0_alu_0_n_40_1), 
      .S(eu_mab[1]), .A(execution_unit_0_n_79), .B(execution_unit_0_alu_0_n_89), 
      .CI(execution_unit_0_alu_0_n_40_0));
  FA_X1_LVT execution_unit_0_alu_0_i_40_2 (.CO(execution_unit_0_alu_0_n_40_2), 
      .S(eu_mab[2]), .A(execution_unit_0_n_80), .B(execution_unit_0_alu_0_n_90), 
      .CI(execution_unit_0_alu_0_n_40_1));
  FA_X1_LVT execution_unit_0_alu_0_i_40_3 (.CO(execution_unit_0_alu_0_n_40_3), 
      .S(eu_mab[3]), .A(execution_unit_0_n_81), .B(execution_unit_0_alu_0_n_91), 
      .CI(execution_unit_0_alu_0_n_40_2));
  FA_X1_LVT execution_unit_0_alu_0_i_40_4 (.CO(execution_unit_0_alu_0_n_40_4), 
      .S(eu_mab[4]), .A(execution_unit_0_n_82), .B(execution_unit_0_alu_0_n_92), 
      .CI(execution_unit_0_alu_0_n_40_3));
  FA_X1_LVT execution_unit_0_alu_0_i_40_5 (.CO(execution_unit_0_alu_0_n_40_5), 
      .S(eu_mab[5]), .A(execution_unit_0_n_83), .B(execution_unit_0_alu_0_n_93), 
      .CI(execution_unit_0_alu_0_n_40_4));
  FA_X1_LVT execution_unit_0_alu_0_i_40_6 (.CO(execution_unit_0_alu_0_n_40_6), 
      .S(eu_mab[6]), .A(execution_unit_0_n_84), .B(execution_unit_0_alu_0_n_94), 
      .CI(execution_unit_0_alu_0_n_40_5));
  FA_X1_LVT execution_unit_0_alu_0_i_40_7 (.CO(execution_unit_0_alu_0_n_40_7), 
      .S(eu_mab[7]), .A(execution_unit_0_n_85), .B(execution_unit_0_alu_0_n_95), 
      .CI(execution_unit_0_alu_0_n_40_6));
  FA_X1_LVT execution_unit_0_alu_0_i_40_8 (.CO(execution_unit_0_alu_0_n_40_8), 
      .S(eu_mab[8]), .A(execution_unit_0_alu_0_n_0), .B(
      execution_unit_0_alu_0_n_96), .CI(execution_unit_0_alu_0_n_40_7));
  FA_X1_LVT execution_unit_0_alu_0_i_40_9 (.CO(execution_unit_0_alu_0_n_40_9), 
      .S(eu_mab[9]), .A(execution_unit_0_alu_0_n_1), .B(
      execution_unit_0_alu_0_n_97), .CI(execution_unit_0_alu_0_n_40_8));
  FA_X1_LVT execution_unit_0_alu_0_i_40_10 (.CO(execution_unit_0_alu_0_n_40_10), 
      .S(eu_mab[10]), .A(execution_unit_0_alu_0_n_2), .B(
      execution_unit_0_alu_0_n_98), .CI(execution_unit_0_alu_0_n_40_9));
  FA_X1_LVT execution_unit_0_alu_0_i_40_11 (.CO(execution_unit_0_alu_0_n_40_11), 
      .S(eu_mab[11]), .A(execution_unit_0_alu_0_n_3), .B(
      execution_unit_0_alu_0_n_99), .CI(execution_unit_0_alu_0_n_40_10));
  FA_X1_LVT execution_unit_0_alu_0_i_40_12 (.CO(execution_unit_0_alu_0_n_40_12), 
      .S(eu_mab[12]), .A(execution_unit_0_alu_0_n_4), .B(
      execution_unit_0_alu_0_n_100), .CI(execution_unit_0_alu_0_n_40_11));
  FA_X1_LVT execution_unit_0_alu_0_i_40_13 (.CO(execution_unit_0_alu_0_n_40_13), 
      .S(eu_mab[13]), .A(execution_unit_0_alu_0_n_5), .B(
      execution_unit_0_alu_0_n_101), .CI(execution_unit_0_alu_0_n_40_12));
  FA_X1_LVT execution_unit_0_alu_0_i_40_14 (.CO(execution_unit_0_alu_0_n_40_14), 
      .S(eu_mab[14]), .A(execution_unit_0_alu_0_n_6), .B(
      execution_unit_0_alu_0_n_102), .CI(execution_unit_0_alu_0_n_40_13));
  FA_X1_LVT execution_unit_0_alu_0_i_40_15 (.CO(
      execution_unit_0_alu_0_alu_add[16]), .S(eu_mab[15]), .A(
      execution_unit_0_alu_0_n_7), .B(execution_unit_0_alu_0_n_103), .CI(
      execution_unit_0_alu_0_n_40_14));
  AOI21_X1_LVT execution_unit_0_alu_0_i_28_0 (.ZN(execution_unit_0_alu_0_n_28_0), 
      .A(inst_alu[1]), .B1(inst_alu[2]), .B2(execution_unit_0_status[0]));
  INV_X1_LVT execution_unit_0_alu_0_i_28_1 (.ZN(execution_unit_0_alu_0_n_28_1), 
      .A(execution_unit_0_n_0));
  NOR2_X1_LVT execution_unit_0_alu_0_i_28_2 (.ZN(execution_unit_0_alu_0_alu_inc), 
      .A1(execution_unit_0_alu_0_n_28_0), .A2(execution_unit_0_alu_0_n_28_1));
  HA_X1_LVT execution_unit_0_alu_0_i_41_0 (.CO(execution_unit_0_alu_0_n_41_0), 
      .S(execution_unit_0_alu_0_alu_add_inc[0]), .A(
      execution_unit_0_alu_0_alu_inc), .B(eu_mab[0]));
  HA_X1_LVT execution_unit_0_alu_0_i_41_1 (.CO(execution_unit_0_alu_0_n_41_1), 
      .S(execution_unit_0_alu_0_alu_add_inc[1]), .A(eu_mab[1]), .B(
      execution_unit_0_alu_0_n_41_0));
  HA_X1_LVT execution_unit_0_alu_0_i_41_2 (.CO(execution_unit_0_alu_0_n_41_2), 
      .S(execution_unit_0_alu_0_alu_add_inc[2]), .A(eu_mab[2]), .B(
      execution_unit_0_alu_0_n_41_1));
  HA_X1_LVT execution_unit_0_alu_0_i_41_3 (.CO(execution_unit_0_alu_0_n_41_3), 
      .S(execution_unit_0_alu_0_alu_add_inc[3]), .A(eu_mab[3]), .B(
      execution_unit_0_alu_0_n_41_2));
  HA_X1_LVT execution_unit_0_alu_0_i_41_4 (.CO(execution_unit_0_alu_0_n_41_4), 
      .S(execution_unit_0_alu_0_alu_add_inc[4]), .A(eu_mab[4]), .B(
      execution_unit_0_alu_0_n_41_3));
  HA_X1_LVT execution_unit_0_alu_0_i_41_5 (.CO(execution_unit_0_alu_0_n_41_5), 
      .S(execution_unit_0_alu_0_alu_add_inc[5]), .A(eu_mab[5]), .B(
      execution_unit_0_alu_0_n_41_4));
  HA_X1_LVT execution_unit_0_alu_0_i_41_6 (.CO(execution_unit_0_alu_0_n_41_6), 
      .S(execution_unit_0_alu_0_alu_add_inc[6]), .A(eu_mab[6]), .B(
      execution_unit_0_alu_0_n_41_5));
  HA_X1_LVT execution_unit_0_alu_0_i_41_7 (.CO(execution_unit_0_alu_0_n_41_7), 
      .S(execution_unit_0_alu_0_alu_add_inc[7]), .A(eu_mab[7]), .B(
      execution_unit_0_alu_0_n_41_6));
  HA_X1_LVT execution_unit_0_alu_0_i_41_8 (.CO(execution_unit_0_alu_0_n_41_8), 
      .S(execution_unit_0_alu_0_alu_add_inc[8]), .A(eu_mab[8]), .B(
      execution_unit_0_alu_0_n_41_7));
  HA_X1_LVT execution_unit_0_alu_0_i_41_9 (.CO(execution_unit_0_alu_0_n_41_9), 
      .S(execution_unit_0_alu_0_alu_add_inc[9]), .A(eu_mab[9]), .B(
      execution_unit_0_alu_0_n_41_8));
  HA_X1_LVT execution_unit_0_alu_0_i_41_10 (.CO(execution_unit_0_alu_0_n_41_10), 
      .S(execution_unit_0_alu_0_alu_add_inc[10]), .A(eu_mab[10]), .B(
      execution_unit_0_alu_0_n_41_9));
  HA_X1_LVT execution_unit_0_alu_0_i_41_11 (.CO(execution_unit_0_alu_0_n_41_11), 
      .S(execution_unit_0_alu_0_alu_add_inc[11]), .A(eu_mab[11]), .B(
      execution_unit_0_alu_0_n_41_10));
  HA_X1_LVT execution_unit_0_alu_0_i_41_12 (.CO(execution_unit_0_alu_0_n_41_12), 
      .S(execution_unit_0_alu_0_alu_add_inc[12]), .A(eu_mab[12]), .B(
      execution_unit_0_alu_0_n_41_11));
  HA_X1_LVT execution_unit_0_alu_0_i_41_13 (.CO(execution_unit_0_alu_0_n_41_13), 
      .S(execution_unit_0_alu_0_alu_add_inc[13]), .A(eu_mab[13]), .B(
      execution_unit_0_alu_0_n_41_12));
  HA_X1_LVT execution_unit_0_alu_0_i_41_14 (.CO(execution_unit_0_alu_0_n_41_14), 
      .S(execution_unit_0_alu_0_alu_add_inc[14]), .A(eu_mab[14]), .B(
      execution_unit_0_alu_0_n_41_13));
  HA_X1_LVT execution_unit_0_alu_0_i_41_15 (.CO(execution_unit_0_alu_0_n_41_15), 
      .S(execution_unit_0_alu_0_alu_add_inc[15]), .A(eu_mab[15]), .B(
      execution_unit_0_alu_0_n_41_14));
  INV_X1_LVT execution_unit_0_alu_0_i_43_1 (.ZN(execution_unit_0_alu_0_n_43_0), 
      .A(inst_alu[7]));
  NOR2_X1_LVT execution_unit_0_alu_0_i_43_2 (.ZN(execution_unit_0_alu_0_n_106), 
      .A1(execution_unit_0_alu_0_n_43_0), .A2(execution_unit_0_alu_0_n_104));
  HA_X1_LVT execution_unit_0_alu_0_i_18_3 (.CO(execution_unit_0_alu_0_n_68), .S(
      execution_unit_0_alu_0_n_67), .A(execution_unit_0_alu_0_n_3), .B(
      execution_unit_0_alu_0_n_19));
  INV_X1_LVT execution_unit_0_alu_0_i_19_2 (.ZN(execution_unit_0_alu_0_n_19_3), 
      .A(execution_unit_0_alu_0_n_68));
  HA_X1_LVT execution_unit_0_alu_0_i_18_2 (.CO(execution_unit_0_alu_0_n_66), .S(
      execution_unit_0_alu_0_n_65), .A(execution_unit_0_alu_0_n_2), .B(
      execution_unit_0_alu_0_n_18));
  HA_X1_LVT execution_unit_0_alu_0_i_19_1 (.CO(execution_unit_0_alu_0_n_19_2), 
      .S(execution_unit_0_alu_0_n_19_1), .A(execution_unit_0_alu_0_n_67), .B(
      execution_unit_0_alu_0_n_66));
  HA_X1_LVT execution_unit_0_alu_0_i_13_3 (.CO(execution_unit_0_alu_0_n_56), .S(
      execution_unit_0_alu_0_n_55), .A(execution_unit_0_n_85), .B(
      execution_unit_0_alu_0_n_15));
  INV_X1_LVT execution_unit_0_alu_0_i_14_2 (.ZN(execution_unit_0_alu_0_n_14_3), 
      .A(execution_unit_0_alu_0_n_56));
  HA_X1_LVT execution_unit_0_alu_0_i_13_2 (.CO(execution_unit_0_alu_0_n_54), .S(
      execution_unit_0_alu_0_n_53), .A(execution_unit_0_n_84), .B(
      execution_unit_0_alu_0_n_14));
  HA_X1_LVT execution_unit_0_alu_0_i_14_1 (.CO(execution_unit_0_alu_0_n_14_2), 
      .S(execution_unit_0_alu_0_n_14_1), .A(execution_unit_0_alu_0_n_55), .B(
      execution_unit_0_alu_0_n_54));
  HA_X1_LVT execution_unit_0_alu_0_i_8_3 (.CO(execution_unit_0_alu_0_n_44), .S(
      execution_unit_0_alu_0_n_43), .A(execution_unit_0_n_81), .B(
      execution_unit_0_alu_0_n_11));
  INV_X1_LVT execution_unit_0_alu_0_i_9_2 (.ZN(execution_unit_0_alu_0_n_9_3), .A(
      execution_unit_0_alu_0_n_44));
  HA_X1_LVT execution_unit_0_alu_0_i_8_2 (.CO(execution_unit_0_alu_0_n_42), .S(
      execution_unit_0_alu_0_n_41), .A(execution_unit_0_n_80), .B(
      execution_unit_0_alu_0_n_10));
  HA_X1_LVT execution_unit_0_alu_0_i_9_1 (.CO(execution_unit_0_alu_0_n_9_2), .S(
      execution_unit_0_alu_0_n_9_1), .A(execution_unit_0_alu_0_n_43), .B(
      execution_unit_0_alu_0_n_42));
  FA_X1_LVT execution_unit_0_alu_0_i_8_0 (.CO(execution_unit_0_alu_0_n_8_0), .S(
      execution_unit_0_alu_0_n_38), .A(execution_unit_0_n_78), .B(
      execution_unit_0_status[0]), .CI(execution_unit_0_alu_0_n_8));
  FA_X1_LVT execution_unit_0_alu_0_i_8_1 (.CO(execution_unit_0_alu_0_n_40), .S(
      execution_unit_0_alu_0_n_39), .A(execution_unit_0_n_79), .B(
      execution_unit_0_alu_0_n_9), .CI(execution_unit_0_alu_0_n_8_0));
  INV_X1_LVT execution_unit_0_alu_0_i_9_0 (.ZN(execution_unit_0_alu_0_n_9_0), .A(
      execution_unit_0_alu_0_n_40));
  FA_X1_LVT execution_unit_0_alu_0_i_9_3 (.CO(execution_unit_0_alu_0_n_9_4), .S(), 
      .A(execution_unit_0_alu_0_n_41), .B(execution_unit_0_alu_0_n_9_0), .CI(
      execution_unit_0_alu_0_n_39));
  FA_X1_LVT execution_unit_0_alu_0_i_9_4 (.CO(execution_unit_0_alu_0_n_9_5), .S(), 
      .A(execution_unit_0_alu_0_n_40), .B(execution_unit_0_alu_0_n_9_1), .CI(
      execution_unit_0_alu_0_n_9_4));
  FA_X1_LVT execution_unit_0_alu_0_i_9_5 (.CO(execution_unit_0_alu_0_n_9_6), .S(), 
      .A(execution_unit_0_alu_0_n_9_2), .B(execution_unit_0_alu_0_n_9_3), .CI(
      execution_unit_0_alu_0_n_9_5));
  HA_X1_LVT execution_unit_0_alu_0_i_9_6 (.CO(execution_unit_0_alu_0_n_9_7), .S(), 
      .A(execution_unit_0_alu_0_n_9_3), .B(execution_unit_0_alu_0_n_9_6));
  HA_X1_LVT execution_unit_0_alu_0_i_9_7 (.CO(execution_unit_0_alu_0_n_9_8), .S(), 
      .A(execution_unit_0_alu_0_n_9_3), .B(execution_unit_0_alu_0_n_9_7));
  XNOR2_X1_LVT execution_unit_0_alu_0_i_9_8 (.ZN(execution_unit_0_alu_0_n_9_9), 
      .A(execution_unit_0_alu_0_n_9_3), .B(execution_unit_0_alu_0_n_9_8));
  INV_X1_LVT execution_unit_0_alu_0_i_9_9 (.ZN(execution_unit_0_alu_0_n_45), .A(
      execution_unit_0_alu_0_n_9_9));
  INV_X1_LVT execution_unit_0_alu_0_i_10_0 (.ZN(execution_unit_0_alu_0_n_46), .A(
      execution_unit_0_alu_0_n_45));
  HA_X1_LVT execution_unit_0_alu_0_i_11_0 (.CO(execution_unit_0_alu_0_n_11_0), 
      .S(execution_unit_0_alu_0_n_47), .A(execution_unit_0_alu_0_n_40), .B(
      execution_unit_0_alu_0_n_41));
  FA_X1_LVT execution_unit_0_alu_0_i_11_1 (.CO(execution_unit_0_alu_0_n_11_1), 
      .S(execution_unit_0_alu_0_n_48), .A(execution_unit_0_alu_0_n_43), .B(
      execution_unit_0_alu_0_n_42), .CI(execution_unit_0_alu_0_n_11_0));
  OR2_X1_LVT execution_unit_0_alu_0_i_12_7 (.ZN(execution_unit_0_alu_0_n_12_5), 
      .A1(execution_unit_0_alu_0_n_46), .A2(execution_unit_0_alu_0_n_48));
  HA_X1_LVT execution_unit_0_alu_0_i_11_2 (.CO(execution_unit_0_alu_0_n_11_2), 
      .S(execution_unit_0_alu_0_n_49), .A(execution_unit_0_alu_0_n_44), .B(
      execution_unit_0_alu_0_n_11_1));
  INV_X1_LVT execution_unit_0_alu_0_i_12_8 (.ZN(execution_unit_0_alu_0_n_12_6), 
      .A(execution_unit_0_alu_0_n_49));
  XNOR2_X1_LVT execution_unit_0_alu_0_i_12_10 (.ZN(execution_unit_0_alu_0_n_12_8), 
      .A(execution_unit_0_alu_0_n_12_5), .B(execution_unit_0_alu_0_n_12_6));
  INV_X1_LVT execution_unit_0_alu_0_i_12_3 (.ZN(execution_unit_0_alu_0_n_12_2), 
      .A(execution_unit_0_alu_0_n_39));
  NAND2_X1_LVT execution_unit_0_alu_0_i_12_2 (.ZN(execution_unit_0_alu_0_n_12_1), 
      .A1(execution_unit_0_alu_0_n_46), .A2(execution_unit_0_alu_0_n_12_2));
  OR2_X1_LVT execution_unit_0_alu_0_i_12_5 (.ZN(execution_unit_0_alu_0_n_12_3), 
      .A1(execution_unit_0_alu_0_n_47), .A2(execution_unit_0_alu_0_n_12_1));
  XNOR2_X1_LVT execution_unit_0_alu_0_i_12_6 (.ZN(execution_unit_0_alu_0_n_12_4), 
      .A(execution_unit_0_alu_0_n_46), .B(execution_unit_0_alu_0_n_48));
  HA_X1_LVT execution_unit_0_alu_0_i_12_9 (.CO(execution_unit_0_alu_0_n_12_7), 
      .S(execution_unit_0_alu_0_bcd_add[3]), .A(execution_unit_0_alu_0_n_12_3), 
      .B(execution_unit_0_alu_0_n_12_4));
  XNOR2_X1_LVT execution_unit_0_alu_0_i_12_11 (.ZN(
      execution_unit_0_alu_0_bcd_add[4]), .A(execution_unit_0_alu_0_n_12_8), .B(
      execution_unit_0_alu_0_n_12_7));
  FA_X1_LVT execution_unit_0_alu_0_i_13_0 (.CO(execution_unit_0_alu_0_n_13_0), 
      .S(execution_unit_0_alu_0_n_50), .A(execution_unit_0_n_82), .B(
      execution_unit_0_alu_0_bcd_add[4]), .CI(execution_unit_0_alu_0_n_12));
  FA_X1_LVT execution_unit_0_alu_0_i_13_1 (.CO(execution_unit_0_alu_0_n_52), .S(
      execution_unit_0_alu_0_n_51), .A(execution_unit_0_n_83), .B(
      execution_unit_0_alu_0_n_13), .CI(execution_unit_0_alu_0_n_13_0));
  INV_X1_LVT execution_unit_0_alu_0_i_14_0 (.ZN(execution_unit_0_alu_0_n_14_0), 
      .A(execution_unit_0_alu_0_n_52));
  FA_X1_LVT execution_unit_0_alu_0_i_14_3 (.CO(execution_unit_0_alu_0_n_14_4), 
      .S(), .A(execution_unit_0_alu_0_n_53), .B(execution_unit_0_alu_0_n_14_0), 
      .CI(execution_unit_0_alu_0_n_51));
  FA_X1_LVT execution_unit_0_alu_0_i_14_4 (.CO(execution_unit_0_alu_0_n_14_5), 
      .S(), .A(execution_unit_0_alu_0_n_52), .B(execution_unit_0_alu_0_n_14_1), 
      .CI(execution_unit_0_alu_0_n_14_4));
  FA_X1_LVT execution_unit_0_alu_0_i_14_5 (.CO(execution_unit_0_alu_0_n_14_6), 
      .S(), .A(execution_unit_0_alu_0_n_14_2), .B(execution_unit_0_alu_0_n_14_3), 
      .CI(execution_unit_0_alu_0_n_14_5));
  HA_X1_LVT execution_unit_0_alu_0_i_14_6 (.CO(execution_unit_0_alu_0_n_14_7), 
      .S(), .A(execution_unit_0_alu_0_n_14_3), .B(execution_unit_0_alu_0_n_14_6));
  HA_X1_LVT execution_unit_0_alu_0_i_14_7 (.CO(execution_unit_0_alu_0_n_14_8), 
      .S(), .A(execution_unit_0_alu_0_n_14_3), .B(execution_unit_0_alu_0_n_14_7));
  XNOR2_X1_LVT execution_unit_0_alu_0_i_14_8 (.ZN(execution_unit_0_alu_0_n_14_9), 
      .A(execution_unit_0_alu_0_n_14_3), .B(execution_unit_0_alu_0_n_14_8));
  INV_X1_LVT execution_unit_0_alu_0_i_14_9 (.ZN(execution_unit_0_alu_0_n_57), .A(
      execution_unit_0_alu_0_n_14_9));
  INV_X1_LVT execution_unit_0_alu_0_i_15_0 (.ZN(execution_unit_0_alu_0_n_58), .A(
      execution_unit_0_alu_0_n_57));
  HA_X1_LVT execution_unit_0_alu_0_i_16_0 (.CO(execution_unit_0_alu_0_n_16_0), 
      .S(execution_unit_0_alu_0_n_59), .A(execution_unit_0_alu_0_n_52), .B(
      execution_unit_0_alu_0_n_53));
  FA_X1_LVT execution_unit_0_alu_0_i_16_1 (.CO(execution_unit_0_alu_0_n_16_1), 
      .S(execution_unit_0_alu_0_n_60), .A(execution_unit_0_alu_0_n_55), .B(
      execution_unit_0_alu_0_n_54), .CI(execution_unit_0_alu_0_n_16_0));
  OR2_X1_LVT execution_unit_0_alu_0_i_17_7 (.ZN(execution_unit_0_alu_0_n_17_5), 
      .A1(execution_unit_0_alu_0_n_58), .A2(execution_unit_0_alu_0_n_60));
  HA_X1_LVT execution_unit_0_alu_0_i_16_2 (.CO(execution_unit_0_alu_0_n_16_2), 
      .S(execution_unit_0_alu_0_n_61), .A(execution_unit_0_alu_0_n_56), .B(
      execution_unit_0_alu_0_n_16_1));
  INV_X1_LVT execution_unit_0_alu_0_i_17_8 (.ZN(execution_unit_0_alu_0_n_17_6), 
      .A(execution_unit_0_alu_0_n_61));
  XNOR2_X1_LVT execution_unit_0_alu_0_i_17_10 (.ZN(execution_unit_0_alu_0_n_17_8), 
      .A(execution_unit_0_alu_0_n_17_5), .B(execution_unit_0_alu_0_n_17_6));
  INV_X1_LVT execution_unit_0_alu_0_i_17_3 (.ZN(execution_unit_0_alu_0_n_17_2), 
      .A(execution_unit_0_alu_0_n_51));
  NAND2_X1_LVT execution_unit_0_alu_0_i_17_2 (.ZN(execution_unit_0_alu_0_n_17_1), 
      .A1(execution_unit_0_alu_0_n_58), .A2(execution_unit_0_alu_0_n_17_2));
  OR2_X1_LVT execution_unit_0_alu_0_i_17_5 (.ZN(execution_unit_0_alu_0_n_17_3), 
      .A1(execution_unit_0_alu_0_n_59), .A2(execution_unit_0_alu_0_n_17_1));
  XNOR2_X1_LVT execution_unit_0_alu_0_i_17_6 (.ZN(execution_unit_0_alu_0_n_17_4), 
      .A(execution_unit_0_alu_0_n_58), .B(execution_unit_0_alu_0_n_60));
  HA_X1_LVT execution_unit_0_alu_0_i_17_9 (.CO(execution_unit_0_alu_0_n_17_7), 
      .S(execution_unit_0_alu_0_bcd_add0[3]), .A(execution_unit_0_alu_0_n_17_3), 
      .B(execution_unit_0_alu_0_n_17_4));
  XNOR2_X1_LVT execution_unit_0_alu_0_i_17_11 (.ZN(
      execution_unit_0_alu_0_bcd_add0[4]), .A(execution_unit_0_alu_0_n_17_8), .B(
      execution_unit_0_alu_0_n_17_7));
  FA_X1_LVT execution_unit_0_alu_0_i_18_0 (.CO(execution_unit_0_alu_0_n_18_0), 
      .S(execution_unit_0_alu_0_n_62), .A(execution_unit_0_alu_0_n_0), .B(
      execution_unit_0_alu_0_bcd_add0[4]), .CI(execution_unit_0_alu_0_n_16));
  FA_X1_LVT execution_unit_0_alu_0_i_18_1 (.CO(execution_unit_0_alu_0_n_64), .S(
      execution_unit_0_alu_0_n_63), .A(execution_unit_0_alu_0_n_1), .B(
      execution_unit_0_alu_0_n_17), .CI(execution_unit_0_alu_0_n_18_0));
  INV_X1_LVT execution_unit_0_alu_0_i_19_0 (.ZN(execution_unit_0_alu_0_n_19_0), 
      .A(execution_unit_0_alu_0_n_64));
  FA_X1_LVT execution_unit_0_alu_0_i_19_3 (.CO(execution_unit_0_alu_0_n_19_4), 
      .S(), .A(execution_unit_0_alu_0_n_65), .B(execution_unit_0_alu_0_n_19_0), 
      .CI(execution_unit_0_alu_0_n_63));
  FA_X1_LVT execution_unit_0_alu_0_i_19_4 (.CO(execution_unit_0_alu_0_n_19_5), 
      .S(), .A(execution_unit_0_alu_0_n_64), .B(execution_unit_0_alu_0_n_19_1), 
      .CI(execution_unit_0_alu_0_n_19_4));
  FA_X1_LVT execution_unit_0_alu_0_i_19_5 (.CO(execution_unit_0_alu_0_n_19_6), 
      .S(), .A(execution_unit_0_alu_0_n_19_2), .B(execution_unit_0_alu_0_n_19_3), 
      .CI(execution_unit_0_alu_0_n_19_5));
  HA_X1_LVT execution_unit_0_alu_0_i_19_6 (.CO(execution_unit_0_alu_0_n_19_7), 
      .S(), .A(execution_unit_0_alu_0_n_19_3), .B(execution_unit_0_alu_0_n_19_6));
  HA_X1_LVT execution_unit_0_alu_0_i_19_7 (.CO(execution_unit_0_alu_0_n_19_8), 
      .S(), .A(execution_unit_0_alu_0_n_19_3), .B(execution_unit_0_alu_0_n_19_7));
  XNOR2_X1_LVT execution_unit_0_alu_0_i_19_8 (.ZN(execution_unit_0_alu_0_n_19_9), 
      .A(execution_unit_0_alu_0_n_19_3), .B(execution_unit_0_alu_0_n_19_8));
  INV_X1_LVT execution_unit_0_alu_0_i_19_9 (.ZN(execution_unit_0_alu_0_n_69), .A(
      execution_unit_0_alu_0_n_19_9));
  INV_X1_LVT execution_unit_0_alu_0_i_20_0 (.ZN(execution_unit_0_alu_0_n_70), .A(
      execution_unit_0_alu_0_n_69));
  HA_X1_LVT execution_unit_0_alu_0_i_21_0 (.CO(execution_unit_0_alu_0_n_21_0), 
      .S(execution_unit_0_alu_0_n_71), .A(execution_unit_0_alu_0_n_64), .B(
      execution_unit_0_alu_0_n_65));
  FA_X1_LVT execution_unit_0_alu_0_i_21_1 (.CO(execution_unit_0_alu_0_n_21_1), 
      .S(execution_unit_0_alu_0_n_72), .A(execution_unit_0_alu_0_n_67), .B(
      execution_unit_0_alu_0_n_66), .CI(execution_unit_0_alu_0_n_21_0));
  OR2_X1_LVT execution_unit_0_alu_0_i_22_7 (.ZN(execution_unit_0_alu_0_n_22_5), 
      .A1(execution_unit_0_alu_0_n_70), .A2(execution_unit_0_alu_0_n_72));
  HA_X1_LVT execution_unit_0_alu_0_i_21_2 (.CO(execution_unit_0_alu_0_n_21_2), 
      .S(execution_unit_0_alu_0_n_73), .A(execution_unit_0_alu_0_n_68), .B(
      execution_unit_0_alu_0_n_21_1));
  INV_X1_LVT execution_unit_0_alu_0_i_22_8 (.ZN(execution_unit_0_alu_0_n_22_6), 
      .A(execution_unit_0_alu_0_n_73));
  XNOR2_X1_LVT execution_unit_0_alu_0_i_22_10 (.ZN(execution_unit_0_alu_0_n_22_8), 
      .A(execution_unit_0_alu_0_n_22_5), .B(execution_unit_0_alu_0_n_22_6));
  INV_X1_LVT execution_unit_0_alu_0_i_22_3 (.ZN(execution_unit_0_alu_0_n_22_2), 
      .A(execution_unit_0_alu_0_n_63));
  NAND2_X1_LVT execution_unit_0_alu_0_i_22_2 (.ZN(execution_unit_0_alu_0_n_22_1), 
      .A1(execution_unit_0_alu_0_n_70), .A2(execution_unit_0_alu_0_n_22_2));
  OR2_X1_LVT execution_unit_0_alu_0_i_22_5 (.ZN(execution_unit_0_alu_0_n_22_3), 
      .A1(execution_unit_0_alu_0_n_71), .A2(execution_unit_0_alu_0_n_22_1));
  XNOR2_X1_LVT execution_unit_0_alu_0_i_22_6 (.ZN(execution_unit_0_alu_0_n_22_4), 
      .A(execution_unit_0_alu_0_n_70), .B(execution_unit_0_alu_0_n_72));
  HA_X1_LVT execution_unit_0_alu_0_i_22_9 (.CO(execution_unit_0_alu_0_n_22_7), 
      .S(execution_unit_0_alu_0_bcd_add1[3]), .A(execution_unit_0_alu_0_n_22_3), 
      .B(execution_unit_0_alu_0_n_22_4));
  XNOR2_X1_LVT execution_unit_0_alu_0_i_22_11 (.ZN(
      execution_unit_0_alu_0_bcd_add1[4]), .A(execution_unit_0_alu_0_n_22_8), .B(
      execution_unit_0_alu_0_n_22_7));
  FA_X1_LVT execution_unit_0_alu_0_i_23_0 (.CO(execution_unit_0_alu_0_n_23_0), 
      .S(execution_unit_0_alu_0_n_74), .A(execution_unit_0_alu_0_n_4), .B(
      execution_unit_0_alu_0_bcd_add1[4]), .CI(execution_unit_0_alu_0_X[0]));
  FA_X1_LVT execution_unit_0_alu_0_i_23_1 (.CO(execution_unit_0_alu_0_n_76), .S(
      execution_unit_0_alu_0_n_75), .A(execution_unit_0_alu_0_n_5), .B(
      execution_unit_0_alu_0_X[1]), .CI(execution_unit_0_alu_0_n_23_0));
  HA_X1_LVT execution_unit_0_alu_0_i_23_2 (.CO(execution_unit_0_alu_0_n_78), .S(
      execution_unit_0_alu_0_n_77), .A(execution_unit_0_alu_0_n_6), .B(
      execution_unit_0_alu_0_X[2]));
  HA_X1_LVT execution_unit_0_alu_0_i_26_0 (.CO(execution_unit_0_alu_0_n_26_0), 
      .S(execution_unit_0_alu_0_n_83), .A(execution_unit_0_alu_0_n_76), .B(
      execution_unit_0_alu_0_n_77));
  HA_X1_LVT execution_unit_0_alu_0_i_23_3 (.CO(execution_unit_0_alu_0_n_80), .S(
      execution_unit_0_alu_0_n_79), .A(execution_unit_0_alu_0_n_7), .B(
      execution_unit_0_alu_0_X[3]));
  INV_X1_LVT execution_unit_0_alu_0_i_24_2 (.ZN(execution_unit_0_alu_0_n_24_3), 
      .A(execution_unit_0_alu_0_n_80));
  HA_X1_LVT execution_unit_0_alu_0_i_24_1 (.CO(execution_unit_0_alu_0_n_24_2), 
      .S(execution_unit_0_alu_0_n_24_1), .A(execution_unit_0_alu_0_n_79), .B(
      execution_unit_0_alu_0_n_78));
  INV_X1_LVT execution_unit_0_alu_0_i_24_0 (.ZN(execution_unit_0_alu_0_n_24_0), 
      .A(execution_unit_0_alu_0_n_76));
  FA_X1_LVT execution_unit_0_alu_0_i_24_3 (.CO(execution_unit_0_alu_0_n_24_4), 
      .S(), .A(execution_unit_0_alu_0_n_77), .B(execution_unit_0_alu_0_n_24_0), 
      .CI(execution_unit_0_alu_0_n_75));
  FA_X1_LVT execution_unit_0_alu_0_i_24_4 (.CO(execution_unit_0_alu_0_n_24_5), 
      .S(), .A(execution_unit_0_alu_0_n_76), .B(execution_unit_0_alu_0_n_24_1), 
      .CI(execution_unit_0_alu_0_n_24_4));
  FA_X1_LVT execution_unit_0_alu_0_i_24_5 (.CO(execution_unit_0_alu_0_n_24_6), 
      .S(), .A(execution_unit_0_alu_0_n_24_2), .B(execution_unit_0_alu_0_n_24_3), 
      .CI(execution_unit_0_alu_0_n_24_5));
  HA_X1_LVT execution_unit_0_alu_0_i_24_6 (.CO(execution_unit_0_alu_0_n_24_7), 
      .S(), .A(execution_unit_0_alu_0_n_24_3), .B(execution_unit_0_alu_0_n_24_6));
  HA_X1_LVT execution_unit_0_alu_0_i_24_7 (.CO(execution_unit_0_alu_0_n_24_8), 
      .S(), .A(execution_unit_0_alu_0_n_24_3), .B(execution_unit_0_alu_0_n_24_7));
  XNOR2_X1_LVT execution_unit_0_alu_0_i_24_8 (.ZN(execution_unit_0_alu_0_n_24_9), 
      .A(execution_unit_0_alu_0_n_24_3), .B(execution_unit_0_alu_0_n_24_8));
  INV_X1_LVT execution_unit_0_alu_0_i_24_9 (.ZN(execution_unit_0_alu_0_n_81), .A(
      execution_unit_0_alu_0_n_24_9));
  INV_X1_LVT execution_unit_0_alu_0_i_25_0 (.ZN(execution_unit_0_alu_0_n_82), .A(
      execution_unit_0_alu_0_n_81));
  INV_X1_LVT execution_unit_0_alu_0_i_27_3 (.ZN(execution_unit_0_alu_0_n_27_2), 
      .A(execution_unit_0_alu_0_n_75));
  NAND2_X1_LVT execution_unit_0_alu_0_i_27_2 (.ZN(execution_unit_0_alu_0_n_27_1), 
      .A1(execution_unit_0_alu_0_n_82), .A2(execution_unit_0_alu_0_n_27_2));
  OR2_X1_LVT execution_unit_0_alu_0_i_27_5 (.ZN(execution_unit_0_alu_0_n_27_3), 
      .A1(execution_unit_0_alu_0_n_83), .A2(execution_unit_0_alu_0_n_27_1));
  FA_X1_LVT execution_unit_0_alu_0_i_26_1 (.CO(execution_unit_0_alu_0_n_26_1), 
      .S(execution_unit_0_alu_0_n_84), .A(execution_unit_0_alu_0_n_79), .B(
      execution_unit_0_alu_0_n_78), .CI(execution_unit_0_alu_0_n_26_0));
  XNOR2_X1_LVT execution_unit_0_alu_0_i_27_6 (.ZN(execution_unit_0_alu_0_n_27_4), 
      .A(execution_unit_0_alu_0_n_82), .B(execution_unit_0_alu_0_n_84));
  HA_X1_LVT execution_unit_0_alu_0_i_27_9 (.CO(execution_unit_0_alu_0_n_27_7), 
      .S(execution_unit_0_alu_0_bcd_add2[3]), .A(execution_unit_0_alu_0_n_27_3), 
      .B(execution_unit_0_alu_0_n_27_4));
  NOR2_X1_LVT execution_unit_0_alu_0_i_43_0 (.ZN(execution_unit_0_alu_0_n_105), 
      .A1(inst_alu[7]), .A2(execution_unit_0_alu_0_n_104));
  OR4_X1_LVT execution_unit_0_alu_0_i_6_0 (.ZN(execution_unit_0_alu_0_n_6_0), 
      .A1(inst_so[1]), .A2(inst_alu[10]), .A3(inst_alu[6]), .A4(inst_alu[5]));
  NOR3_X1_LVT execution_unit_0_alu_0_i_6_1 (.ZN(
      execution_unit_0_alu_0_alu_short_thro), .A1(execution_unit_0_alu_0_n_6_0), 
      .A2(inst_alu[4]), .A3(inst_so[3]));
  NAND2_X1_LVT execution_unit_0_alu_0_i_7_143 (.ZN(
      execution_unit_0_alu_0_n_7_128), .A1(execution_unit_0_alu_0_alu_short_thro), 
      .A2(execution_unit_0_alu_0_X[3]));
  NAND2_X1_LVT execution_unit_0_alu_0_i_7_71 (.ZN(execution_unit_0_alu_0_n_7_64), 
      .A1(inst_so[3]), .A2(execution_unit_0_n_116));
  NAND2_X1_LVT execution_unit_0_alu_0_i_7_144 (.ZN(
      execution_unit_0_alu_0_n_7_129), .A1(inst_so[1]), .A2(
      execution_unit_0_n_116));
  INV_X1_LVT execution_unit_0_alu_0_i_5_0 (.ZN(execution_unit_0_alu_0_n_5_0), .A(
      inst_bw));
  INV_X1_LVT execution_unit_0_alu_0_i_5_1 (.ZN(execution_unit_0_alu_0_n_5_1), .A(
      inst_so[0]));
  NAND3_X1_LVT execution_unit_0_alu_0_i_5_2 (.ZN(execution_unit_0_alu_0_n_5_2), 
      .A1(execution_unit_0_alu_0_n_5_0), .A2(execution_unit_0_alu_0_n_5_1), .A3(
      execution_unit_0_n_124));
  NAND3_X1_LVT execution_unit_0_alu_0_i_5_3 (.ZN(execution_unit_0_alu_0_n_5_3), 
      .A1(execution_unit_0_alu_0_n_5_1), .A2(inst_bw), .A3(
      execution_unit_0_n_116));
  NAND2_X1_LVT execution_unit_0_alu_0_i_5_4 (.ZN(execution_unit_0_alu_0_n_5_4), 
      .A1(execution_unit_0_status[0]), .A2(inst_so[0]));
  NAND3_X1_LVT execution_unit_0_alu_0_i_5_5 (.ZN(execution_unit_0_alu_0_n_20), 
      .A1(execution_unit_0_alu_0_n_5_2), .A2(execution_unit_0_alu_0_n_5_3), .A3(
      execution_unit_0_alu_0_n_5_4));
  NAND2_X1_LVT execution_unit_0_alu_0_i_7_145 (.ZN(
      execution_unit_0_alu_0_n_7_130), .A1(inst_alu[10]), .A2(
      execution_unit_0_alu_0_n_20));
  AND4_X1_LVT execution_unit_0_alu_0_i_7_146 (.ZN(execution_unit_0_alu_0_n_7_131), 
      .A1(execution_unit_0_alu_0_n_7_128), .A2(execution_unit_0_alu_0_n_7_64), 
      .A3(execution_unit_0_alu_0_n_7_129), .A4(execution_unit_0_alu_0_n_7_130));
  OAI21_X1_LVT execution_unit_0_alu_0_i_7_147 (.ZN(
      execution_unit_0_alu_0_n_7_132), .A(inst_alu[5]), .B1(
      execution_unit_0_alu_0_X[3]), .B2(execution_unit_0_alu_0_n_7));
  XOR2_X1_LVT execution_unit_0_alu_0_i_7_148 (.Z(execution_unit_0_alu_0_n_7_133), 
      .A(execution_unit_0_alu_0_X[3]), .B(execution_unit_0_alu_0_n_7));
  NAND2_X1_LVT execution_unit_0_alu_0_i_7_149 (.ZN(
      execution_unit_0_alu_0_n_7_134), .A1(execution_unit_0_alu_0_n_7_133), .A2(
      inst_alu[6]));
  NAND3_X1_LVT execution_unit_0_alu_0_i_7_150 (.ZN(
      execution_unit_0_alu_0_n_7_135), .A1(inst_alu[4]), .A2(
      execution_unit_0_alu_0_X[3]), .A3(execution_unit_0_alu_0_n_7));
  NAND4_X1_LVT execution_unit_0_alu_0_i_7_151 (.ZN(execution_unit_0_alu_0_n_37), 
      .A1(execution_unit_0_alu_0_n_7_131), .A2(execution_unit_0_alu_0_n_7_132), 
      .A3(execution_unit_0_alu_0_n_7_134), .A4(execution_unit_0_alu_0_n_7_135));
  AOI222_X1_LVT execution_unit_0_alu_0_i_44_30 (.ZN(
      execution_unit_0_alu_0_n_44_15), .A1(execution_unit_0_alu_0_n_104), .A2(
      execution_unit_0_alu_0_alu_add_inc[15]), .B1(execution_unit_0_alu_0_n_106), 
      .B2(execution_unit_0_alu_0_bcd_add2[3]), .C1(execution_unit_0_alu_0_n_105), 
      .C2(execution_unit_0_alu_0_n_37));
  INV_X1_LVT execution_unit_0_alu_0_i_44_31 (.ZN(execution_unit_0_alu_out[15]), 
      .A(execution_unit_0_alu_0_n_44_15));
  XNOR2_X1_LVT execution_unit_0_alu_0_i_27_4 (.ZN(
      execution_unit_0_alu_0_bcd_add2[2]), .A(execution_unit_0_alu_0_n_83), .B(
      execution_unit_0_alu_0_n_27_1));
  NAND2_X1_LVT execution_unit_0_alu_0_i_7_134 (.ZN(
      execution_unit_0_alu_0_n_7_120), .A1(execution_unit_0_alu_0_alu_short_thro), 
      .A2(execution_unit_0_alu_0_X[2]));
  NAND2_X1_LVT execution_unit_0_alu_0_i_7_135 (.ZN(
      execution_unit_0_alu_0_n_7_121), .A1(inst_so[1]), .A2(
      execution_unit_0_n_115));
  NAND2_X1_LVT execution_unit_0_alu_0_i_7_136 (.ZN(
      execution_unit_0_alu_0_n_7_122), .A1(inst_alu[10]), .A2(
      execution_unit_0_n_124));
  AND4_X1_LVT execution_unit_0_alu_0_i_7_137 (.ZN(execution_unit_0_alu_0_n_7_123), 
      .A1(execution_unit_0_alu_0_n_7_120), .A2(execution_unit_0_alu_0_n_7_64), 
      .A3(execution_unit_0_alu_0_n_7_121), .A4(execution_unit_0_alu_0_n_7_122));
  OAI21_X1_LVT execution_unit_0_alu_0_i_7_138 (.ZN(
      execution_unit_0_alu_0_n_7_124), .A(inst_alu[5]), .B1(
      execution_unit_0_alu_0_X[2]), .B2(execution_unit_0_alu_0_n_6));
  XOR2_X1_LVT execution_unit_0_alu_0_i_7_139 (.Z(execution_unit_0_alu_0_n_7_125), 
      .A(execution_unit_0_alu_0_X[2]), .B(execution_unit_0_alu_0_n_6));
  NAND2_X1_LVT execution_unit_0_alu_0_i_7_140 (.ZN(
      execution_unit_0_alu_0_n_7_126), .A1(execution_unit_0_alu_0_n_7_125), .A2(
      inst_alu[6]));
  NAND3_X1_LVT execution_unit_0_alu_0_i_7_141 (.ZN(
      execution_unit_0_alu_0_n_7_127), .A1(inst_alu[4]), .A2(
      execution_unit_0_alu_0_X[2]), .A3(execution_unit_0_alu_0_n_6));
  NAND4_X1_LVT execution_unit_0_alu_0_i_7_142 (.ZN(execution_unit_0_alu_0_n_36), 
      .A1(execution_unit_0_alu_0_n_7_123), .A2(execution_unit_0_alu_0_n_7_124), 
      .A3(execution_unit_0_alu_0_n_7_126), .A4(execution_unit_0_alu_0_n_7_127));
  AOI222_X1_LVT execution_unit_0_alu_0_i_44_28 (.ZN(
      execution_unit_0_alu_0_n_44_14), .A1(execution_unit_0_alu_0_n_104), .A2(
      execution_unit_0_alu_0_alu_add_inc[14]), .B1(execution_unit_0_alu_0_n_106), 
      .B2(execution_unit_0_alu_0_bcd_add2[2]), .C1(execution_unit_0_alu_0_n_105), 
      .C2(execution_unit_0_alu_0_n_36));
  INV_X1_LVT execution_unit_0_alu_0_i_44_29 (.ZN(execution_unit_0_alu_out[14]), 
      .A(execution_unit_0_alu_0_n_44_14));
  XNOR2_X1_LVT execution_unit_0_alu_0_i_27_0 (.ZN(execution_unit_0_alu_0_n_27_0), 
      .A(execution_unit_0_alu_0_n_82), .B(execution_unit_0_alu_0_n_75));
  INV_X1_LVT execution_unit_0_alu_0_i_27_1 (.ZN(
      execution_unit_0_alu_0_bcd_add2[1]), .A(execution_unit_0_alu_0_n_27_0));
  NAND2_X1_LVT execution_unit_0_alu_0_i_7_125 (.ZN(
      execution_unit_0_alu_0_n_7_112), .A1(execution_unit_0_alu_0_alu_short_thro), 
      .A2(execution_unit_0_alu_0_X[1]));
  NAND2_X1_LVT execution_unit_0_alu_0_i_7_126 (.ZN(
      execution_unit_0_alu_0_n_7_113), .A1(inst_so[1]), .A2(
      execution_unit_0_n_114));
  NAND2_X1_LVT execution_unit_0_alu_0_i_7_127 (.ZN(
      execution_unit_0_alu_0_n_7_114), .A1(inst_alu[10]), .A2(
      execution_unit_0_n_123));
  AND4_X1_LVT execution_unit_0_alu_0_i_7_128 (.ZN(execution_unit_0_alu_0_n_7_115), 
      .A1(execution_unit_0_alu_0_n_7_112), .A2(execution_unit_0_alu_0_n_7_64), 
      .A3(execution_unit_0_alu_0_n_7_113), .A4(execution_unit_0_alu_0_n_7_114));
  OAI21_X1_LVT execution_unit_0_alu_0_i_7_129 (.ZN(
      execution_unit_0_alu_0_n_7_116), .A(inst_alu[5]), .B1(
      execution_unit_0_alu_0_X[1]), .B2(execution_unit_0_alu_0_n_5));
  XOR2_X1_LVT execution_unit_0_alu_0_i_7_130 (.Z(execution_unit_0_alu_0_n_7_117), 
      .A(execution_unit_0_alu_0_X[1]), .B(execution_unit_0_alu_0_n_5));
  NAND2_X1_LVT execution_unit_0_alu_0_i_7_131 (.ZN(
      execution_unit_0_alu_0_n_7_118), .A1(execution_unit_0_alu_0_n_7_117), .A2(
      inst_alu[6]));
  NAND3_X1_LVT execution_unit_0_alu_0_i_7_132 (.ZN(
      execution_unit_0_alu_0_n_7_119), .A1(inst_alu[4]), .A2(
      execution_unit_0_alu_0_X[1]), .A3(execution_unit_0_alu_0_n_5));
  NAND4_X1_LVT execution_unit_0_alu_0_i_7_133 (.ZN(execution_unit_0_alu_0_n_35), 
      .A1(execution_unit_0_alu_0_n_7_115), .A2(execution_unit_0_alu_0_n_7_116), 
      .A3(execution_unit_0_alu_0_n_7_118), .A4(execution_unit_0_alu_0_n_7_119));
  AOI222_X1_LVT execution_unit_0_alu_0_i_44_26 (.ZN(
      execution_unit_0_alu_0_n_44_13), .A1(execution_unit_0_alu_0_n_104), .A2(
      execution_unit_0_alu_0_alu_add_inc[13]), .B1(execution_unit_0_alu_0_n_106), 
      .B2(execution_unit_0_alu_0_bcd_add2[1]), .C1(execution_unit_0_alu_0_n_105), 
      .C2(execution_unit_0_alu_0_n_35));
  INV_X1_LVT execution_unit_0_alu_0_i_44_27 (.ZN(execution_unit_0_alu_out[13]), 
      .A(execution_unit_0_alu_0_n_44_13));
  NAND2_X1_LVT execution_unit_0_alu_0_i_7_116 (.ZN(
      execution_unit_0_alu_0_n_7_104), .A1(execution_unit_0_alu_0_alu_short_thro), 
      .A2(execution_unit_0_alu_0_X[0]));
  NAND2_X1_LVT execution_unit_0_alu_0_i_7_117 (.ZN(
      execution_unit_0_alu_0_n_7_105), .A1(inst_so[1]), .A2(
      execution_unit_0_n_113));
  NAND2_X1_LVT execution_unit_0_alu_0_i_7_118 (.ZN(
      execution_unit_0_alu_0_n_7_106), .A1(inst_alu[10]), .A2(
      execution_unit_0_n_122));
  AND4_X1_LVT execution_unit_0_alu_0_i_7_119 (.ZN(execution_unit_0_alu_0_n_7_107), 
      .A1(execution_unit_0_alu_0_n_7_104), .A2(execution_unit_0_alu_0_n_7_64), 
      .A3(execution_unit_0_alu_0_n_7_105), .A4(execution_unit_0_alu_0_n_7_106));
  OAI21_X1_LVT execution_unit_0_alu_0_i_7_120 (.ZN(
      execution_unit_0_alu_0_n_7_108), .A(inst_alu[5]), .B1(
      execution_unit_0_alu_0_X[0]), .B2(execution_unit_0_alu_0_n_4));
  XOR2_X1_LVT execution_unit_0_alu_0_i_7_121 (.Z(execution_unit_0_alu_0_n_7_109), 
      .A(execution_unit_0_alu_0_X[0]), .B(execution_unit_0_alu_0_n_4));
  NAND2_X1_LVT execution_unit_0_alu_0_i_7_122 (.ZN(
      execution_unit_0_alu_0_n_7_110), .A1(execution_unit_0_alu_0_n_7_109), .A2(
      inst_alu[6]));
  NAND3_X1_LVT execution_unit_0_alu_0_i_7_123 (.ZN(
      execution_unit_0_alu_0_n_7_111), .A1(inst_alu[4]), .A2(
      execution_unit_0_alu_0_X[0]), .A3(execution_unit_0_alu_0_n_4));
  NAND4_X1_LVT execution_unit_0_alu_0_i_7_124 (.ZN(execution_unit_0_alu_0_n_34), 
      .A1(execution_unit_0_alu_0_n_7_107), .A2(execution_unit_0_alu_0_n_7_108), 
      .A3(execution_unit_0_alu_0_n_7_110), .A4(execution_unit_0_alu_0_n_7_111));
  AOI222_X1_LVT execution_unit_0_alu_0_i_44_24 (.ZN(
      execution_unit_0_alu_0_n_44_12), .A1(execution_unit_0_alu_0_n_104), .A2(
      execution_unit_0_alu_0_alu_add_inc[12]), .B1(execution_unit_0_alu_0_n_106), 
      .B2(execution_unit_0_alu_0_n_74), .C1(execution_unit_0_alu_0_n_105), .C2(
      execution_unit_0_alu_0_n_34));
  INV_X1_LVT execution_unit_0_alu_0_i_44_25 (.ZN(execution_unit_0_alu_out[12]), 
      .A(execution_unit_0_alu_0_n_44_12));
  NAND2_X1_LVT execution_unit_0_alu_0_i_7_107 (.ZN(execution_unit_0_alu_0_n_7_96), 
      .A1(execution_unit_0_alu_0_alu_short_thro), .A2(
      execution_unit_0_alu_0_n_19));
  NAND2_X1_LVT execution_unit_0_alu_0_i_7_108 (.ZN(execution_unit_0_alu_0_n_7_97), 
      .A1(inst_so[1]), .A2(execution_unit_0_n_112));
  NAND2_X1_LVT execution_unit_0_alu_0_i_7_109 (.ZN(execution_unit_0_alu_0_n_7_98), 
      .A1(inst_alu[10]), .A2(execution_unit_0_n_121));
  AND4_X1_LVT execution_unit_0_alu_0_i_7_110 (.ZN(execution_unit_0_alu_0_n_7_99), 
      .A1(execution_unit_0_alu_0_n_7_96), .A2(execution_unit_0_alu_0_n_7_64), 
      .A3(execution_unit_0_alu_0_n_7_97), .A4(execution_unit_0_alu_0_n_7_98));
  OAI21_X1_LVT execution_unit_0_alu_0_i_7_111 (.ZN(
      execution_unit_0_alu_0_n_7_100), .A(inst_alu[5]), .B1(
      execution_unit_0_alu_0_n_19), .B2(execution_unit_0_alu_0_n_3));
  XOR2_X1_LVT execution_unit_0_alu_0_i_7_112 (.Z(execution_unit_0_alu_0_n_7_101), 
      .A(execution_unit_0_alu_0_n_19), .B(execution_unit_0_alu_0_n_3));
  NAND2_X1_LVT execution_unit_0_alu_0_i_7_113 (.ZN(
      execution_unit_0_alu_0_n_7_102), .A1(execution_unit_0_alu_0_n_7_101), .A2(
      inst_alu[6]));
  NAND3_X1_LVT execution_unit_0_alu_0_i_7_114 (.ZN(
      execution_unit_0_alu_0_n_7_103), .A1(inst_alu[4]), .A2(
      execution_unit_0_alu_0_n_19), .A3(execution_unit_0_alu_0_n_3));
  NAND4_X1_LVT execution_unit_0_alu_0_i_7_115 (.ZN(execution_unit_0_alu_0_n_33), 
      .A1(execution_unit_0_alu_0_n_7_99), .A2(execution_unit_0_alu_0_n_7_100), 
      .A3(execution_unit_0_alu_0_n_7_102), .A4(execution_unit_0_alu_0_n_7_103));
  AOI222_X1_LVT execution_unit_0_alu_0_i_44_22 (.ZN(
      execution_unit_0_alu_0_n_44_11), .A1(execution_unit_0_alu_0_n_104), .A2(
      execution_unit_0_alu_0_alu_add_inc[11]), .B1(execution_unit_0_alu_0_n_106), 
      .B2(execution_unit_0_alu_0_bcd_add1[3]), .C1(execution_unit_0_alu_0_n_105), 
      .C2(execution_unit_0_alu_0_n_33));
  INV_X1_LVT execution_unit_0_alu_0_i_44_23 (.ZN(execution_unit_0_alu_out[11]), 
      .A(execution_unit_0_alu_0_n_44_11));
  XNOR2_X1_LVT execution_unit_0_alu_0_i_22_4 (.ZN(
      execution_unit_0_alu_0_bcd_add1[2]), .A(execution_unit_0_alu_0_n_71), .B(
      execution_unit_0_alu_0_n_22_1));
  NAND2_X1_LVT execution_unit_0_alu_0_i_7_98 (.ZN(execution_unit_0_alu_0_n_7_88), 
      .A1(execution_unit_0_alu_0_alu_short_thro), .A2(
      execution_unit_0_alu_0_n_18));
  NAND2_X1_LVT execution_unit_0_alu_0_i_7_99 (.ZN(execution_unit_0_alu_0_n_7_89), 
      .A1(inst_so[1]), .A2(execution_unit_0_n_111));
  NAND2_X1_LVT execution_unit_0_alu_0_i_7_100 (.ZN(execution_unit_0_alu_0_n_7_90), 
      .A1(inst_alu[10]), .A2(execution_unit_0_n_120));
  AND4_X1_LVT execution_unit_0_alu_0_i_7_101 (.ZN(execution_unit_0_alu_0_n_7_91), 
      .A1(execution_unit_0_alu_0_n_7_88), .A2(execution_unit_0_alu_0_n_7_64), 
      .A3(execution_unit_0_alu_0_n_7_89), .A4(execution_unit_0_alu_0_n_7_90));
  OAI21_X1_LVT execution_unit_0_alu_0_i_7_102 (.ZN(execution_unit_0_alu_0_n_7_92), 
      .A(inst_alu[5]), .B1(execution_unit_0_alu_0_n_18), .B2(
      execution_unit_0_alu_0_n_2));
  XOR2_X1_LVT execution_unit_0_alu_0_i_7_103 (.Z(execution_unit_0_alu_0_n_7_93), 
      .A(execution_unit_0_alu_0_n_18), .B(execution_unit_0_alu_0_n_2));
  NAND2_X1_LVT execution_unit_0_alu_0_i_7_104 (.ZN(execution_unit_0_alu_0_n_7_94), 
      .A1(execution_unit_0_alu_0_n_7_93), .A2(inst_alu[6]));
  NAND3_X1_LVT execution_unit_0_alu_0_i_7_105 (.ZN(execution_unit_0_alu_0_n_7_95), 
      .A1(inst_alu[4]), .A2(execution_unit_0_alu_0_n_18), .A3(
      execution_unit_0_alu_0_n_2));
  NAND4_X1_LVT execution_unit_0_alu_0_i_7_106 (.ZN(execution_unit_0_alu_0_n_32), 
      .A1(execution_unit_0_alu_0_n_7_91), .A2(execution_unit_0_alu_0_n_7_92), 
      .A3(execution_unit_0_alu_0_n_7_94), .A4(execution_unit_0_alu_0_n_7_95));
  AOI222_X1_LVT execution_unit_0_alu_0_i_44_20 (.ZN(
      execution_unit_0_alu_0_n_44_10), .A1(execution_unit_0_alu_0_n_104), .A2(
      execution_unit_0_alu_0_alu_add_inc[10]), .B1(execution_unit_0_alu_0_n_106), 
      .B2(execution_unit_0_alu_0_bcd_add1[2]), .C1(execution_unit_0_alu_0_n_105), 
      .C2(execution_unit_0_alu_0_n_32));
  INV_X1_LVT execution_unit_0_alu_0_i_44_21 (.ZN(execution_unit_0_alu_out[10]), 
      .A(execution_unit_0_alu_0_n_44_10));
  XNOR2_X1_LVT execution_unit_0_alu_0_i_22_0 (.ZN(execution_unit_0_alu_0_n_22_0), 
      .A(execution_unit_0_alu_0_n_70), .B(execution_unit_0_alu_0_n_63));
  INV_X1_LVT execution_unit_0_alu_0_i_22_1 (.ZN(
      execution_unit_0_alu_0_bcd_add1[1]), .A(execution_unit_0_alu_0_n_22_0));
  NAND2_X1_LVT execution_unit_0_alu_0_i_7_89 (.ZN(execution_unit_0_alu_0_n_7_80), 
      .A1(execution_unit_0_alu_0_alu_short_thro), .A2(
      execution_unit_0_alu_0_n_17));
  NAND2_X1_LVT execution_unit_0_alu_0_i_7_90 (.ZN(execution_unit_0_alu_0_n_7_81), 
      .A1(inst_so[1]), .A2(execution_unit_0_n_110));
  NAND2_X1_LVT execution_unit_0_alu_0_i_7_91 (.ZN(execution_unit_0_alu_0_n_7_82), 
      .A1(inst_alu[10]), .A2(execution_unit_0_n_119));
  AND4_X1_LVT execution_unit_0_alu_0_i_7_92 (.ZN(execution_unit_0_alu_0_n_7_83), 
      .A1(execution_unit_0_alu_0_n_7_80), .A2(execution_unit_0_alu_0_n_7_64), 
      .A3(execution_unit_0_alu_0_n_7_81), .A4(execution_unit_0_alu_0_n_7_82));
  OAI21_X1_LVT execution_unit_0_alu_0_i_7_93 (.ZN(execution_unit_0_alu_0_n_7_84), 
      .A(inst_alu[5]), .B1(execution_unit_0_alu_0_n_17), .B2(
      execution_unit_0_alu_0_n_1));
  XOR2_X1_LVT execution_unit_0_alu_0_i_7_94 (.Z(execution_unit_0_alu_0_n_7_85), 
      .A(execution_unit_0_alu_0_n_17), .B(execution_unit_0_alu_0_n_1));
  NAND2_X1_LVT execution_unit_0_alu_0_i_7_95 (.ZN(execution_unit_0_alu_0_n_7_86), 
      .A1(execution_unit_0_alu_0_n_7_85), .A2(inst_alu[6]));
  NAND3_X1_LVT execution_unit_0_alu_0_i_7_96 (.ZN(execution_unit_0_alu_0_n_7_87), 
      .A1(inst_alu[4]), .A2(execution_unit_0_alu_0_n_17), .A3(
      execution_unit_0_alu_0_n_1));
  NAND4_X1_LVT execution_unit_0_alu_0_i_7_97 (.ZN(execution_unit_0_alu_0_n_31), 
      .A1(execution_unit_0_alu_0_n_7_83), .A2(execution_unit_0_alu_0_n_7_84), 
      .A3(execution_unit_0_alu_0_n_7_86), .A4(execution_unit_0_alu_0_n_7_87));
  AOI222_X1_LVT execution_unit_0_alu_0_i_44_18 (.ZN(
      execution_unit_0_alu_0_n_44_9), .A1(execution_unit_0_alu_0_n_104), .A2(
      execution_unit_0_alu_0_alu_add_inc[9]), .B1(execution_unit_0_alu_0_n_106), 
      .B2(execution_unit_0_alu_0_bcd_add1[1]), .C1(execution_unit_0_alu_0_n_105), 
      .C2(execution_unit_0_alu_0_n_31));
  INV_X1_LVT execution_unit_0_alu_0_i_44_19 (.ZN(execution_unit_0_alu_out[9]), 
      .A(execution_unit_0_alu_0_n_44_9));
  NAND2_X1_LVT execution_unit_0_alu_0_i_7_80 (.ZN(execution_unit_0_alu_0_n_7_72), 
      .A1(execution_unit_0_alu_0_alu_short_thro), .A2(
      execution_unit_0_alu_0_n_16));
  NAND2_X1_LVT execution_unit_0_alu_0_i_7_81 (.ZN(execution_unit_0_alu_0_n_7_73), 
      .A1(execution_unit_0_n_109), .A2(inst_so[1]));
  NAND2_X1_LVT execution_unit_0_alu_0_i_7_82 (.ZN(execution_unit_0_alu_0_n_7_74), 
      .A1(inst_alu[10]), .A2(execution_unit_0_n_118));
  AND4_X1_LVT execution_unit_0_alu_0_i_7_83 (.ZN(execution_unit_0_alu_0_n_7_75), 
      .A1(execution_unit_0_alu_0_n_7_72), .A2(execution_unit_0_alu_0_n_7_64), 
      .A3(execution_unit_0_alu_0_n_7_73), .A4(execution_unit_0_alu_0_n_7_74));
  OAI21_X1_LVT execution_unit_0_alu_0_i_7_84 (.ZN(execution_unit_0_alu_0_n_7_76), 
      .A(inst_alu[5]), .B1(execution_unit_0_alu_0_n_16), .B2(
      execution_unit_0_alu_0_n_0));
  XOR2_X1_LVT execution_unit_0_alu_0_i_7_85 (.Z(execution_unit_0_alu_0_n_7_77), 
      .A(execution_unit_0_alu_0_n_16), .B(execution_unit_0_alu_0_n_0));
  NAND2_X1_LVT execution_unit_0_alu_0_i_7_86 (.ZN(execution_unit_0_alu_0_n_7_78), 
      .A1(execution_unit_0_alu_0_n_7_77), .A2(inst_alu[6]));
  NAND3_X1_LVT execution_unit_0_alu_0_i_7_87 (.ZN(execution_unit_0_alu_0_n_7_79), 
      .A1(inst_alu[4]), .A2(execution_unit_0_alu_0_n_16), .A3(
      execution_unit_0_alu_0_n_0));
  NAND4_X1_LVT execution_unit_0_alu_0_i_7_88 (.ZN(execution_unit_0_alu_0_n_30), 
      .A1(execution_unit_0_alu_0_n_7_75), .A2(execution_unit_0_alu_0_n_7_76), 
      .A3(execution_unit_0_alu_0_n_7_78), .A4(execution_unit_0_alu_0_n_7_79));
  AOI222_X1_LVT execution_unit_0_alu_0_i_44_16 (.ZN(
      execution_unit_0_alu_0_n_44_8), .A1(execution_unit_0_alu_0_n_104), .A2(
      execution_unit_0_alu_0_alu_add_inc[8]), .B1(execution_unit_0_alu_0_n_106), 
      .B2(execution_unit_0_alu_0_n_62), .C1(execution_unit_0_alu_0_n_105), .C2(
      execution_unit_0_alu_0_n_30));
  INV_X1_LVT execution_unit_0_alu_0_i_44_17 (.ZN(execution_unit_0_alu_out[8]), 
      .A(execution_unit_0_alu_0_n_44_8));
  NAND2_X1_LVT execution_unit_0_alu_0_i_7_70 (.ZN(execution_unit_0_alu_0_n_7_63), 
      .A1(execution_unit_0_alu_0_alu_short_thro), .A2(
      execution_unit_0_alu_0_n_15));
  NAND2_X1_LVT execution_unit_0_alu_0_i_7_72 (.ZN(execution_unit_0_alu_0_n_7_65), 
      .A1(inst_so[1]), .A2(execution_unit_0_n_124));
  AOI22_X1_LVT execution_unit_0_alu_0_i_5_6 (.ZN(execution_unit_0_alu_0_n_5_5), 
      .A1(execution_unit_0_alu_0_n_20), .A2(inst_bw), .B1(
      execution_unit_0_alu_0_n_5_0), .B2(execution_unit_0_n_117));
  INV_X1_LVT execution_unit_0_alu_0_i_5_7 (.ZN(execution_unit_0_alu_0_n_21), .A(
      execution_unit_0_alu_0_n_5_5));
  NAND2_X1_LVT execution_unit_0_alu_0_i_7_73 (.ZN(execution_unit_0_alu_0_n_7_66), 
      .A1(inst_alu[10]), .A2(execution_unit_0_alu_0_n_21));
  AND4_X1_LVT execution_unit_0_alu_0_i_7_74 (.ZN(execution_unit_0_alu_0_n_7_67), 
      .A1(execution_unit_0_alu_0_n_7_63), .A2(execution_unit_0_alu_0_n_7_64), 
      .A3(execution_unit_0_alu_0_n_7_65), .A4(execution_unit_0_alu_0_n_7_66));
  OAI21_X1_LVT execution_unit_0_alu_0_i_7_75 (.ZN(execution_unit_0_alu_0_n_7_68), 
      .A(inst_alu[5]), .B1(execution_unit_0_alu_0_n_15), .B2(
      execution_unit_0_n_85));
  XOR2_X1_LVT execution_unit_0_alu_0_i_7_76 (.Z(execution_unit_0_alu_0_n_7_69), 
      .A(execution_unit_0_alu_0_n_15), .B(execution_unit_0_n_85));
  NAND2_X1_LVT execution_unit_0_alu_0_i_7_77 (.ZN(execution_unit_0_alu_0_n_7_70), 
      .A1(execution_unit_0_alu_0_n_7_69), .A2(inst_alu[6]));
  NAND3_X1_LVT execution_unit_0_alu_0_i_7_78 (.ZN(execution_unit_0_alu_0_n_7_71), 
      .A1(inst_alu[4]), .A2(execution_unit_0_alu_0_n_15), .A3(
      execution_unit_0_n_85));
  NAND4_X1_LVT execution_unit_0_alu_0_i_7_79 (.ZN(execution_unit_0_alu_0_n_29), 
      .A1(execution_unit_0_alu_0_n_7_67), .A2(execution_unit_0_alu_0_n_7_68), 
      .A3(execution_unit_0_alu_0_n_7_70), .A4(execution_unit_0_alu_0_n_7_71));
  AOI222_X1_LVT execution_unit_0_alu_0_i_44_14 (.ZN(
      execution_unit_0_alu_0_n_44_7), .A1(execution_unit_0_alu_0_n_104), .A2(
      execution_unit_0_alu_0_alu_add_inc[7]), .B1(execution_unit_0_alu_0_n_106), 
      .B2(execution_unit_0_alu_0_bcd_add0[3]), .C1(execution_unit_0_alu_0_n_105), 
      .C2(execution_unit_0_alu_0_n_29));
  INV_X1_LVT execution_unit_0_alu_0_i_44_15 (.ZN(execution_unit_0_alu_out[7]), 
      .A(execution_unit_0_alu_0_n_44_7));
  XNOR2_X1_LVT execution_unit_0_alu_0_i_17_4 (.ZN(
      execution_unit_0_alu_0_bcd_add0[2]), .A(execution_unit_0_alu_0_n_59), .B(
      execution_unit_0_alu_0_n_17_1));
  NAND2_X1_LVT execution_unit_0_alu_0_i_7_60 (.ZN(execution_unit_0_alu_0_n_7_54), 
      .A1(execution_unit_0_alu_0_alu_short_thro), .A2(
      execution_unit_0_alu_0_n_14));
  NAND2_X1_LVT execution_unit_0_alu_0_i_7_61 (.ZN(execution_unit_0_alu_0_n_7_55), 
      .A1(inst_so[3]), .A2(execution_unit_0_n_115));
  NAND2_X1_LVT execution_unit_0_alu_0_i_7_62 (.ZN(execution_unit_0_alu_0_n_7_56), 
      .A1(inst_so[1]), .A2(execution_unit_0_n_123));
  NAND2_X1_LVT execution_unit_0_alu_0_i_7_63 (.ZN(execution_unit_0_alu_0_n_7_57), 
      .A1(inst_alu[10]), .A2(execution_unit_0_n_116));
  AND4_X1_LVT execution_unit_0_alu_0_i_7_64 (.ZN(execution_unit_0_alu_0_n_7_58), 
      .A1(execution_unit_0_alu_0_n_7_54), .A2(execution_unit_0_alu_0_n_7_55), 
      .A3(execution_unit_0_alu_0_n_7_56), .A4(execution_unit_0_alu_0_n_7_57));
  OAI21_X1_LVT execution_unit_0_alu_0_i_7_65 (.ZN(execution_unit_0_alu_0_n_7_59), 
      .A(inst_alu[5]), .B1(execution_unit_0_alu_0_n_14), .B2(
      execution_unit_0_n_84));
  XOR2_X1_LVT execution_unit_0_alu_0_i_7_66 (.Z(execution_unit_0_alu_0_n_7_60), 
      .A(execution_unit_0_alu_0_n_14), .B(execution_unit_0_n_84));
  NAND2_X1_LVT execution_unit_0_alu_0_i_7_67 (.ZN(execution_unit_0_alu_0_n_7_61), 
      .A1(execution_unit_0_alu_0_n_7_60), .A2(inst_alu[6]));
  NAND3_X1_LVT execution_unit_0_alu_0_i_7_68 (.ZN(execution_unit_0_alu_0_n_7_62), 
      .A1(inst_alu[4]), .A2(execution_unit_0_alu_0_n_14), .A3(
      execution_unit_0_n_84));
  NAND4_X1_LVT execution_unit_0_alu_0_i_7_69 (.ZN(execution_unit_0_alu_0_n_28), 
      .A1(execution_unit_0_alu_0_n_7_58), .A2(execution_unit_0_alu_0_n_7_59), 
      .A3(execution_unit_0_alu_0_n_7_61), .A4(execution_unit_0_alu_0_n_7_62));
  AOI222_X1_LVT execution_unit_0_alu_0_i_44_12 (.ZN(
      execution_unit_0_alu_0_n_44_6), .A1(execution_unit_0_alu_0_n_104), .A2(
      execution_unit_0_alu_0_alu_add_inc[6]), .B1(execution_unit_0_alu_0_n_106), 
      .B2(execution_unit_0_alu_0_bcd_add0[2]), .C1(execution_unit_0_alu_0_n_105), 
      .C2(execution_unit_0_alu_0_n_28));
  INV_X1_LVT execution_unit_0_alu_0_i_44_13 (.ZN(execution_unit_0_alu_out[6]), 
      .A(execution_unit_0_alu_0_n_44_6));
  XNOR2_X1_LVT execution_unit_0_alu_0_i_17_0 (.ZN(execution_unit_0_alu_0_n_17_0), 
      .A(execution_unit_0_alu_0_n_58), .B(execution_unit_0_alu_0_n_51));
  INV_X1_LVT execution_unit_0_alu_0_i_17_1 (.ZN(
      execution_unit_0_alu_0_bcd_add0[1]), .A(execution_unit_0_alu_0_n_17_0));
  NAND2_X1_LVT execution_unit_0_alu_0_i_7_50 (.ZN(execution_unit_0_alu_0_n_7_45), 
      .A1(execution_unit_0_alu_0_alu_short_thro), .A2(
      execution_unit_0_alu_0_n_13));
  NAND2_X1_LVT execution_unit_0_alu_0_i_7_51 (.ZN(execution_unit_0_alu_0_n_7_46), 
      .A1(inst_so[3]), .A2(execution_unit_0_n_114));
  NAND2_X1_LVT execution_unit_0_alu_0_i_7_52 (.ZN(execution_unit_0_alu_0_n_7_47), 
      .A1(inst_so[1]), .A2(execution_unit_0_n_122));
  NAND2_X1_LVT execution_unit_0_alu_0_i_7_53 (.ZN(execution_unit_0_alu_0_n_7_48), 
      .A1(inst_alu[10]), .A2(execution_unit_0_n_115));
  AND4_X1_LVT execution_unit_0_alu_0_i_7_54 (.ZN(execution_unit_0_alu_0_n_7_49), 
      .A1(execution_unit_0_alu_0_n_7_45), .A2(execution_unit_0_alu_0_n_7_46), 
      .A3(execution_unit_0_alu_0_n_7_47), .A4(execution_unit_0_alu_0_n_7_48));
  OAI21_X1_LVT execution_unit_0_alu_0_i_7_55 (.ZN(execution_unit_0_alu_0_n_7_50), 
      .A(inst_alu[5]), .B1(execution_unit_0_alu_0_n_13), .B2(
      execution_unit_0_n_83));
  XOR2_X1_LVT execution_unit_0_alu_0_i_7_56 (.Z(execution_unit_0_alu_0_n_7_51), 
      .A(execution_unit_0_alu_0_n_13), .B(execution_unit_0_n_83));
  NAND2_X1_LVT execution_unit_0_alu_0_i_7_57 (.ZN(execution_unit_0_alu_0_n_7_52), 
      .A1(execution_unit_0_alu_0_n_7_51), .A2(inst_alu[6]));
  NAND3_X1_LVT execution_unit_0_alu_0_i_7_58 (.ZN(execution_unit_0_alu_0_n_7_53), 
      .A1(inst_alu[4]), .A2(execution_unit_0_alu_0_n_13), .A3(
      execution_unit_0_n_83));
  NAND4_X1_LVT execution_unit_0_alu_0_i_7_59 (.ZN(execution_unit_0_alu_0_n_27), 
      .A1(execution_unit_0_alu_0_n_7_49), .A2(execution_unit_0_alu_0_n_7_50), 
      .A3(execution_unit_0_alu_0_n_7_52), .A4(execution_unit_0_alu_0_n_7_53));
  AOI222_X1_LVT execution_unit_0_alu_0_i_44_10 (.ZN(
      execution_unit_0_alu_0_n_44_5), .A1(execution_unit_0_alu_0_n_104), .A2(
      execution_unit_0_alu_0_alu_add_inc[5]), .B1(execution_unit_0_alu_0_n_106), 
      .B2(execution_unit_0_alu_0_bcd_add0[1]), .C1(execution_unit_0_alu_0_n_105), 
      .C2(execution_unit_0_alu_0_n_27));
  INV_X1_LVT execution_unit_0_alu_0_i_44_11 (.ZN(execution_unit_0_alu_out[5]), 
      .A(execution_unit_0_alu_0_n_44_5));
  NAND2_X1_LVT execution_unit_0_alu_0_i_7_40 (.ZN(execution_unit_0_alu_0_n_7_36), 
      .A1(execution_unit_0_alu_0_alu_short_thro), .A2(
      execution_unit_0_alu_0_n_12));
  NAND2_X1_LVT execution_unit_0_alu_0_i_7_41 (.ZN(execution_unit_0_alu_0_n_7_37), 
      .A1(inst_so[3]), .A2(execution_unit_0_n_113));
  NAND2_X1_LVT execution_unit_0_alu_0_i_7_42 (.ZN(execution_unit_0_alu_0_n_7_38), 
      .A1(inst_so[1]), .A2(execution_unit_0_n_121));
  NAND2_X1_LVT execution_unit_0_alu_0_i_7_43 (.ZN(execution_unit_0_alu_0_n_7_39), 
      .A1(inst_alu[10]), .A2(execution_unit_0_n_114));
  AND4_X1_LVT execution_unit_0_alu_0_i_7_44 (.ZN(execution_unit_0_alu_0_n_7_40), 
      .A1(execution_unit_0_alu_0_n_7_36), .A2(execution_unit_0_alu_0_n_7_37), 
      .A3(execution_unit_0_alu_0_n_7_38), .A4(execution_unit_0_alu_0_n_7_39));
  OAI21_X1_LVT execution_unit_0_alu_0_i_7_45 (.ZN(execution_unit_0_alu_0_n_7_41), 
      .A(inst_alu[5]), .B1(execution_unit_0_alu_0_n_12), .B2(
      execution_unit_0_n_82));
  XOR2_X1_LVT execution_unit_0_alu_0_i_7_46 (.Z(execution_unit_0_alu_0_n_7_42), 
      .A(execution_unit_0_alu_0_n_12), .B(execution_unit_0_n_82));
  NAND2_X1_LVT execution_unit_0_alu_0_i_7_47 (.ZN(execution_unit_0_alu_0_n_7_43), 
      .A1(execution_unit_0_alu_0_n_7_42), .A2(inst_alu[6]));
  NAND3_X1_LVT execution_unit_0_alu_0_i_7_48 (.ZN(execution_unit_0_alu_0_n_7_44), 
      .A1(inst_alu[4]), .A2(execution_unit_0_alu_0_n_12), .A3(
      execution_unit_0_n_82));
  NAND4_X1_LVT execution_unit_0_alu_0_i_7_49 (.ZN(execution_unit_0_alu_0_n_26), 
      .A1(execution_unit_0_alu_0_n_7_40), .A2(execution_unit_0_alu_0_n_7_41), 
      .A3(execution_unit_0_alu_0_n_7_43), .A4(execution_unit_0_alu_0_n_7_44));
  AOI222_X1_LVT execution_unit_0_alu_0_i_44_8 (.ZN(execution_unit_0_alu_0_n_44_4), 
      .A1(execution_unit_0_alu_0_n_104), .A2(
      execution_unit_0_alu_0_alu_add_inc[4]), .B1(execution_unit_0_alu_0_n_106), 
      .B2(execution_unit_0_alu_0_n_50), .C1(execution_unit_0_alu_0_n_105), .C2(
      execution_unit_0_alu_0_n_26));
  INV_X1_LVT execution_unit_0_alu_0_i_44_9 (.ZN(execution_unit_0_alu_out[4]), .A(
      execution_unit_0_alu_0_n_44_4));
  NAND2_X1_LVT execution_unit_0_alu_0_i_7_30 (.ZN(execution_unit_0_alu_0_n_7_27), 
      .A1(execution_unit_0_alu_0_alu_short_thro), .A2(
      execution_unit_0_alu_0_n_11));
  NAND2_X1_LVT execution_unit_0_alu_0_i_7_31 (.ZN(execution_unit_0_alu_0_n_7_28), 
      .A1(inst_so[3]), .A2(execution_unit_0_n_112));
  NAND2_X1_LVT execution_unit_0_alu_0_i_7_32 (.ZN(execution_unit_0_alu_0_n_7_29), 
      .A1(inst_so[1]), .A2(execution_unit_0_n_120));
  NAND2_X1_LVT execution_unit_0_alu_0_i_7_33 (.ZN(execution_unit_0_alu_0_n_7_30), 
      .A1(inst_alu[10]), .A2(execution_unit_0_n_113));
  AND4_X1_LVT execution_unit_0_alu_0_i_7_34 (.ZN(execution_unit_0_alu_0_n_7_31), 
      .A1(execution_unit_0_alu_0_n_7_27), .A2(execution_unit_0_alu_0_n_7_28), 
      .A3(execution_unit_0_alu_0_n_7_29), .A4(execution_unit_0_alu_0_n_7_30));
  OAI21_X1_LVT execution_unit_0_alu_0_i_7_35 (.ZN(execution_unit_0_alu_0_n_7_32), 
      .A(inst_alu[5]), .B1(execution_unit_0_alu_0_n_11), .B2(
      execution_unit_0_n_81));
  XOR2_X1_LVT execution_unit_0_alu_0_i_7_36 (.Z(execution_unit_0_alu_0_n_7_33), 
      .A(execution_unit_0_alu_0_n_11), .B(execution_unit_0_n_81));
  NAND2_X1_LVT execution_unit_0_alu_0_i_7_37 (.ZN(execution_unit_0_alu_0_n_7_34), 
      .A1(execution_unit_0_alu_0_n_7_33), .A2(inst_alu[6]));
  NAND3_X1_LVT execution_unit_0_alu_0_i_7_38 (.ZN(execution_unit_0_alu_0_n_7_35), 
      .A1(inst_alu[4]), .A2(execution_unit_0_alu_0_n_11), .A3(
      execution_unit_0_n_81));
  NAND4_X1_LVT execution_unit_0_alu_0_i_7_39 (.ZN(execution_unit_0_alu_0_n_25), 
      .A1(execution_unit_0_alu_0_n_7_31), .A2(execution_unit_0_alu_0_n_7_32), 
      .A3(execution_unit_0_alu_0_n_7_34), .A4(execution_unit_0_alu_0_n_7_35));
  AOI222_X1_LVT execution_unit_0_alu_0_i_44_6 (.ZN(execution_unit_0_alu_0_n_44_3), 
      .A1(execution_unit_0_alu_0_n_104), .A2(
      execution_unit_0_alu_0_alu_add_inc[3]), .B1(execution_unit_0_alu_0_n_106), 
      .B2(execution_unit_0_alu_0_bcd_add[3]), .C1(execution_unit_0_alu_0_n_105), 
      .C2(execution_unit_0_alu_0_n_25));
  INV_X1_LVT execution_unit_0_alu_0_i_44_7 (.ZN(execution_unit_0_alu_out[3]), .A(
      execution_unit_0_alu_0_n_44_3));
  XNOR2_X1_LVT execution_unit_0_alu_0_i_12_4 (.ZN(
      execution_unit_0_alu_0_bcd_add[2]), .A(execution_unit_0_alu_0_n_47), .B(
      execution_unit_0_alu_0_n_12_1));
  NAND2_X1_LVT execution_unit_0_alu_0_i_7_20 (.ZN(execution_unit_0_alu_0_n_7_18), 
      .A1(execution_unit_0_alu_0_alu_short_thro), .A2(
      execution_unit_0_alu_0_n_10));
  NAND2_X1_LVT execution_unit_0_alu_0_i_7_21 (.ZN(execution_unit_0_alu_0_n_7_19), 
      .A1(inst_so[3]), .A2(execution_unit_0_n_111));
  NAND2_X1_LVT execution_unit_0_alu_0_i_7_22 (.ZN(execution_unit_0_alu_0_n_7_20), 
      .A1(inst_so[1]), .A2(execution_unit_0_n_119));
  NAND2_X1_LVT execution_unit_0_alu_0_i_7_23 (.ZN(execution_unit_0_alu_0_n_7_21), 
      .A1(inst_alu[10]), .A2(execution_unit_0_n_112));
  AND4_X1_LVT execution_unit_0_alu_0_i_7_24 (.ZN(execution_unit_0_alu_0_n_7_22), 
      .A1(execution_unit_0_alu_0_n_7_18), .A2(execution_unit_0_alu_0_n_7_19), 
      .A3(execution_unit_0_alu_0_n_7_20), .A4(execution_unit_0_alu_0_n_7_21));
  OAI21_X1_LVT execution_unit_0_alu_0_i_7_25 (.ZN(execution_unit_0_alu_0_n_7_23), 
      .A(inst_alu[5]), .B1(execution_unit_0_alu_0_n_10), .B2(
      execution_unit_0_n_80));
  XOR2_X1_LVT execution_unit_0_alu_0_i_7_26 (.Z(execution_unit_0_alu_0_n_7_24), 
      .A(execution_unit_0_alu_0_n_10), .B(execution_unit_0_n_80));
  NAND2_X1_LVT execution_unit_0_alu_0_i_7_27 (.ZN(execution_unit_0_alu_0_n_7_25), 
      .A1(execution_unit_0_alu_0_n_7_24), .A2(inst_alu[6]));
  NAND3_X1_LVT execution_unit_0_alu_0_i_7_28 (.ZN(execution_unit_0_alu_0_n_7_26), 
      .A1(inst_alu[4]), .A2(execution_unit_0_alu_0_n_10), .A3(
      execution_unit_0_n_80));
  NAND4_X1_LVT execution_unit_0_alu_0_i_7_29 (.ZN(execution_unit_0_alu_0_n_24), 
      .A1(execution_unit_0_alu_0_n_7_22), .A2(execution_unit_0_alu_0_n_7_23), 
      .A3(execution_unit_0_alu_0_n_7_25), .A4(execution_unit_0_alu_0_n_7_26));
  AOI222_X1_LVT execution_unit_0_alu_0_i_44_4 (.ZN(execution_unit_0_alu_0_n_44_2), 
      .A1(execution_unit_0_alu_0_n_104), .A2(
      execution_unit_0_alu_0_alu_add_inc[2]), .B1(execution_unit_0_alu_0_n_106), 
      .B2(execution_unit_0_alu_0_bcd_add[2]), .C1(execution_unit_0_alu_0_n_105), 
      .C2(execution_unit_0_alu_0_n_24));
  INV_X1_LVT execution_unit_0_alu_0_i_44_5 (.ZN(execution_unit_0_alu_out[2]), .A(
      execution_unit_0_alu_0_n_44_2));
  XNOR2_X1_LVT execution_unit_0_alu_0_i_12_0 (.ZN(execution_unit_0_alu_0_n_12_0), 
      .A(execution_unit_0_alu_0_n_46), .B(execution_unit_0_alu_0_n_39));
  INV_X1_LVT execution_unit_0_alu_0_i_12_1 (.ZN(
      execution_unit_0_alu_0_bcd_add[1]), .A(execution_unit_0_alu_0_n_12_0));
  NAND2_X1_LVT execution_unit_0_alu_0_i_7_10 (.ZN(execution_unit_0_alu_0_n_7_9), 
      .A1(execution_unit_0_alu_0_alu_short_thro), .A2(execution_unit_0_alu_0_n_9));
  NAND2_X1_LVT execution_unit_0_alu_0_i_7_11 (.ZN(execution_unit_0_alu_0_n_7_10), 
      .A1(inst_so[3]), .A2(execution_unit_0_n_110));
  NAND2_X1_LVT execution_unit_0_alu_0_i_7_12 (.ZN(execution_unit_0_alu_0_n_7_11), 
      .A1(inst_so[1]), .A2(execution_unit_0_n_118));
  NAND2_X1_LVT execution_unit_0_alu_0_i_7_13 (.ZN(execution_unit_0_alu_0_n_7_12), 
      .A1(inst_alu[10]), .A2(execution_unit_0_n_111));
  AND4_X1_LVT execution_unit_0_alu_0_i_7_14 (.ZN(execution_unit_0_alu_0_n_7_13), 
      .A1(execution_unit_0_alu_0_n_7_9), .A2(execution_unit_0_alu_0_n_7_10), .A3(
      execution_unit_0_alu_0_n_7_11), .A4(execution_unit_0_alu_0_n_7_12));
  OAI21_X1_LVT execution_unit_0_alu_0_i_7_15 (.ZN(execution_unit_0_alu_0_n_7_14), 
      .A(inst_alu[5]), .B1(execution_unit_0_alu_0_n_9), .B2(
      execution_unit_0_n_79));
  XOR2_X1_LVT execution_unit_0_alu_0_i_7_16 (.Z(execution_unit_0_alu_0_n_7_15), 
      .A(execution_unit_0_alu_0_n_9), .B(execution_unit_0_n_79));
  NAND2_X1_LVT execution_unit_0_alu_0_i_7_17 (.ZN(execution_unit_0_alu_0_n_7_16), 
      .A1(execution_unit_0_alu_0_n_7_15), .A2(inst_alu[6]));
  NAND3_X1_LVT execution_unit_0_alu_0_i_7_18 (.ZN(execution_unit_0_alu_0_n_7_17), 
      .A1(inst_alu[4]), .A2(execution_unit_0_alu_0_n_9), .A3(
      execution_unit_0_n_79));
  NAND4_X1_LVT execution_unit_0_alu_0_i_7_19 (.ZN(execution_unit_0_alu_0_n_23), 
      .A1(execution_unit_0_alu_0_n_7_13), .A2(execution_unit_0_alu_0_n_7_14), 
      .A3(execution_unit_0_alu_0_n_7_16), .A4(execution_unit_0_alu_0_n_7_17));
  AOI222_X1_LVT execution_unit_0_alu_0_i_44_2 (.ZN(execution_unit_0_alu_0_n_44_1), 
      .A1(execution_unit_0_alu_0_n_104), .A2(
      execution_unit_0_alu_0_alu_add_inc[1]), .B1(execution_unit_0_alu_0_n_106), 
      .B2(execution_unit_0_alu_0_bcd_add[1]), .C1(execution_unit_0_alu_0_n_105), 
      .C2(execution_unit_0_alu_0_n_23));
  INV_X1_LVT execution_unit_0_alu_0_i_44_3 (.ZN(execution_unit_0_alu_out[1]), .A(
      execution_unit_0_alu_0_n_44_1));
  NAND2_X1_LVT execution_unit_0_alu_0_i_7_0 (.ZN(execution_unit_0_alu_0_n_7_0), 
      .A1(execution_unit_0_alu_0_n_8), .A2(execution_unit_0_alu_0_alu_short_thro));
  NAND2_X1_LVT execution_unit_0_alu_0_i_7_1 (.ZN(execution_unit_0_alu_0_n_7_1), 
      .A1(inst_so[3]), .A2(execution_unit_0_n_109));
  NAND2_X1_LVT execution_unit_0_alu_0_i_7_2 (.ZN(execution_unit_0_alu_0_n_7_2), 
      .A1(inst_so[1]), .A2(execution_unit_0_n_117));
  NAND2_X1_LVT execution_unit_0_alu_0_i_7_3 (.ZN(execution_unit_0_alu_0_n_7_3), 
      .A1(inst_alu[10]), .A2(execution_unit_0_n_110));
  AND4_X1_LVT execution_unit_0_alu_0_i_7_4 (.ZN(execution_unit_0_alu_0_n_7_4), 
      .A1(execution_unit_0_alu_0_n_7_0), .A2(execution_unit_0_alu_0_n_7_1), .A3(
      execution_unit_0_alu_0_n_7_2), .A4(execution_unit_0_alu_0_n_7_3));
  OAI21_X1_LVT execution_unit_0_alu_0_i_7_5 (.ZN(execution_unit_0_alu_0_n_7_5), 
      .A(inst_alu[5]), .B1(execution_unit_0_alu_0_n_8), .B2(
      execution_unit_0_n_78));
  XOR2_X1_LVT execution_unit_0_alu_0_i_7_6 (.Z(execution_unit_0_alu_0_n_7_6), .A(
      execution_unit_0_alu_0_n_8), .B(execution_unit_0_n_78));
  NAND2_X1_LVT execution_unit_0_alu_0_i_7_7 (.ZN(execution_unit_0_alu_0_n_7_7), 
      .A1(execution_unit_0_alu_0_n_7_6), .A2(inst_alu[6]));
  NAND3_X1_LVT execution_unit_0_alu_0_i_7_8 (.ZN(execution_unit_0_alu_0_n_7_8), 
      .A1(inst_alu[4]), .A2(execution_unit_0_alu_0_n_8), .A3(
      execution_unit_0_n_78));
  NAND4_X1_LVT execution_unit_0_alu_0_i_7_9 (.ZN(execution_unit_0_alu_0_n_22), 
      .A1(execution_unit_0_alu_0_n_7_4), .A2(execution_unit_0_alu_0_n_7_5), .A3(
      execution_unit_0_alu_0_n_7_7), .A4(execution_unit_0_alu_0_n_7_8));
  AOI222_X1_LVT execution_unit_0_alu_0_i_44_0 (.ZN(execution_unit_0_alu_0_n_44_0), 
      .A1(execution_unit_0_alu_0_alu_add_inc[0]), .A2(
      execution_unit_0_alu_0_n_104), .B1(execution_unit_0_alu_0_n_38), .B2(
      execution_unit_0_alu_0_n_106), .C1(execution_unit_0_alu_0_n_22), .C2(
      execution_unit_0_alu_0_n_105));
  INV_X1_LVT execution_unit_0_alu_0_i_44_1 (.ZN(execution_unit_0_alu_out[0]), .A(
      execution_unit_0_alu_0_n_44_0));
  NOR2_X1_LVT execution_unit_0_alu_0_i_51_1 (.ZN(execution_unit_0_alu_0_n_51_1), 
      .A1(inst_alu[8]), .A2(inst_alu[10]));
  NAND2_X1_LVT execution_unit_0_alu_0_i_51_2 (.ZN(execution_unit_0_alu_0_n_51_2), 
      .A1(execution_unit_0_alu_0_n_51_1), .A2(inst_alu[6]));
  INV_X1_LVT execution_unit_0_alu_0_i_51_8 (.ZN(execution_unit_0_alu_0_n_51_8), 
      .A(inst_bw));
  AND2_X1_LVT execution_unit_0_alu_0_i_45_0 (.ZN(execution_unit_0_alu_0_n_108), 
      .A1(execution_unit_0_alu_0_X[3]), .A2(execution_unit_0_alu_0_n_7));
  AND2_X1_LVT execution_unit_0_alu_0_i_47_0 (.ZN(execution_unit_0_alu_0_n_110), 
      .A1(execution_unit_0_alu_0_n_15), .A2(execution_unit_0_n_85));
  AOI22_X1_LVT execution_unit_0_alu_0_i_51_24 (.ZN(
      execution_unit_0_alu_0_n_51_21), .A1(execution_unit_0_alu_0_n_51_8), .A2(
      execution_unit_0_alu_0_n_108), .B1(inst_bw), .B2(
      execution_unit_0_alu_0_n_110));
  INV_X1_LVT execution_unit_0_alu_0_i_51_6 (.ZN(execution_unit_0_alu_0_n_51_6), 
      .A(inst_alu[6]));
  NAND2_X1_LVT execution_unit_0_alu_0_i_51_7 (.ZN(execution_unit_0_alu_0_n_51_7), 
      .A1(execution_unit_0_alu_0_n_51_1), .A2(execution_unit_0_alu_0_n_51_6));
  INV_X1_LVT execution_unit_0_alu_0_i_46_0 (.ZN(execution_unit_0_alu_0_n_46_0), 
      .A(execution_unit_0_alu_out[15]));
  NOR3_X1_LVT execution_unit_0_alu_0_i_46_1 (.ZN(execution_unit_0_alu_0_n_46_1), 
      .A1(execution_unit_0_alu_0_n_46_0), .A2(execution_unit_0_alu_0_X[3]), .A3(
      execution_unit_0_alu_0_n_7));
  AOI21_X1_LVT execution_unit_0_alu_0_i_46_2 (.ZN(execution_unit_0_alu_0_n_46_2), 
      .A(execution_unit_0_alu_0_n_46_1), .B1(execution_unit_0_alu_0_n_46_0), .B2(
      execution_unit_0_alu_0_n_108));
  INV_X1_LVT execution_unit_0_alu_0_i_46_3 (.ZN(execution_unit_0_alu_0_n_109), 
      .A(execution_unit_0_alu_0_n_46_2));
  INV_X1_LVT execution_unit_0_alu_0_i_48_0 (.ZN(execution_unit_0_alu_0_n_48_0), 
      .A(execution_unit_0_alu_out[7]));
  NOR3_X1_LVT execution_unit_0_alu_0_i_48_1 (.ZN(execution_unit_0_alu_0_n_48_1), 
      .A1(execution_unit_0_alu_0_n_48_0), .A2(execution_unit_0_alu_0_n_15), .A3(
      execution_unit_0_n_85));
  AOI21_X1_LVT execution_unit_0_alu_0_i_48_2 (.ZN(execution_unit_0_alu_0_n_48_2), 
      .A(execution_unit_0_alu_0_n_48_1), .B1(execution_unit_0_alu_0_n_48_0), .B2(
      execution_unit_0_alu_0_n_110));
  INV_X1_LVT execution_unit_0_alu_0_i_48_3 (.ZN(execution_unit_0_alu_0_n_111), 
      .A(execution_unit_0_alu_0_n_48_2));
  AOI22_X1_LVT execution_unit_0_alu_0_i_51_25 (.ZN(
      execution_unit_0_alu_0_n_51_22), .A1(execution_unit_0_alu_0_n_51_8), .A2(
      execution_unit_0_alu_0_n_109), .B1(inst_bw), .B2(
      execution_unit_0_alu_0_n_111));
  OAI22_X1_LVT execution_unit_0_alu_0_i_51_26 (.ZN(execution_unit_0_alu_stat[3]), 
      .A1(execution_unit_0_alu_0_n_51_2), .A2(execution_unit_0_alu_0_n_51_21), 
      .B1(execution_unit_0_alu_0_n_51_7), .B2(execution_unit_0_alu_0_n_51_22));
  INV_X1_LVT execution_unit_0_alu_0_i_51_21 (.ZN(execution_unit_0_alu_0_n_51_19), 
      .A(execution_unit_0_alu_out[7]));
  INV_X1_LVT execution_unit_0_alu_0_i_51_22 (.ZN(execution_unit_0_alu_0_n_51_20), 
      .A(execution_unit_0_alu_out[15]));
  OAI22_X1_LVT execution_unit_0_alu_0_i_51_23 (.ZN(execution_unit_0_alu_stat[2]), 
      .A1(execution_unit_0_alu_0_n_51_8), .A2(execution_unit_0_alu_0_n_51_19), 
      .B1(execution_unit_0_alu_0_n_51_20), .B2(inst_bw));
  OR4_X1_LVT execution_unit_0_alu_0_i_51_11 (.ZN(execution_unit_0_alu_0_n_51_10), 
      .A1(execution_unit_0_alu_0_n_51_8), .A2(execution_unit_0_alu_out[5]), .A3(
      execution_unit_0_alu_out[6]), .A4(execution_unit_0_alu_out[7]));
  OR4_X1_LVT execution_unit_0_alu_0_i_51_12 (.ZN(execution_unit_0_alu_0_n_51_11), 
      .A1(execution_unit_0_alu_0_n_51_10), .A2(execution_unit_0_alu_out[2]), .A3(
      execution_unit_0_alu_out[3]), .A4(execution_unit_0_alu_out[4]));
  OR3_X1_LVT execution_unit_0_alu_0_i_51_13 (.ZN(execution_unit_0_alu_0_n_51_12), 
      .A1(execution_unit_0_alu_0_n_51_11), .A2(execution_unit_0_alu_out[0]), .A3(
      execution_unit_0_alu_out[1]));
  NOR4_X1_LVT execution_unit_0_alu_0_i_51_14 (.ZN(execution_unit_0_alu_0_n_51_13), 
      .A1(execution_unit_0_alu_out[13]), .A2(execution_unit_0_alu_out[14]), .A3(
      execution_unit_0_alu_out[15]), .A4(inst_bw));
  NOR4_X1_LVT execution_unit_0_alu_0_i_51_15 (.ZN(execution_unit_0_alu_0_n_51_14), 
      .A1(execution_unit_0_alu_out[4]), .A2(execution_unit_0_alu_out[5]), .A3(
      execution_unit_0_alu_out[6]), .A4(execution_unit_0_alu_out[7]));
  NOR4_X1_LVT execution_unit_0_alu_0_i_51_16 (.ZN(execution_unit_0_alu_0_n_51_15), 
      .A1(execution_unit_0_alu_out[9]), .A2(execution_unit_0_alu_out[10]), .A3(
      execution_unit_0_alu_out[11]), .A4(execution_unit_0_alu_out[12]));
  INV_X1_LVT execution_unit_0_alu_0_i_51_17 (.ZN(execution_unit_0_alu_0_n_51_16), 
      .A(execution_unit_0_alu_out[3]));
  NAND4_X1_LVT execution_unit_0_alu_0_i_51_18 (.ZN(
      execution_unit_0_alu_0_n_51_17), .A1(execution_unit_0_alu_0_n_51_13), .A2(
      execution_unit_0_alu_0_n_51_14), .A3(execution_unit_0_alu_0_n_51_15), .A4(
      execution_unit_0_alu_0_n_51_16));
  OR4_X1_LVT execution_unit_0_alu_0_i_51_19 (.ZN(execution_unit_0_alu_0_n_51_18), 
      .A1(execution_unit_0_alu_0_n_51_17), .A2(execution_unit_0_alu_out[0]), .A3(
      execution_unit_0_alu_out[1]), .A4(execution_unit_0_alu_out[2]));
  OAI21_X1_LVT execution_unit_0_alu_0_i_51_20 (.ZN(execution_unit_0_alu_stat[1]), 
      .A(execution_unit_0_alu_0_n_51_12), .B1(execution_unit_0_alu_0_n_51_18), 
      .B2(execution_unit_0_alu_out[8]));
  NAND2_X1_LVT execution_unit_0_alu_0_i_51_0 (.ZN(execution_unit_0_alu_0_n_51_0), 
      .A1(execution_unit_0_alu_0_n_8), .A2(inst_alu[10]));
  INV_X1_LVT execution_unit_0_alu_0_i_51_3 (.ZN(execution_unit_0_alu_0_n_51_3), 
      .A(inst_alu[8]));
  OAI21_X1_LVT execution_unit_0_alu_0_i_51_4 (.ZN(execution_unit_0_alu_0_n_51_4), 
      .A(execution_unit_0_alu_0_n_51_2), .B1(inst_alu[10]), .B2(
      execution_unit_0_alu_0_n_51_3));
  INV_X1_LVT execution_unit_0_alu_0_i_49_0 (.ZN(execution_unit_0_alu_0_n_49_0), 
      .A(inst_bw));
  OR4_X1_LVT execution_unit_0_alu_0_i_49_1 (.ZN(execution_unit_0_alu_0_n_49_1), 
      .A1(execution_unit_0_alu_0_n_49_0), .A2(execution_unit_0_alu_out[5]), .A3(
      execution_unit_0_alu_out[6]), .A4(execution_unit_0_alu_out[7]));
  OR4_X1_LVT execution_unit_0_alu_0_i_49_2 (.ZN(execution_unit_0_alu_0_n_49_2), 
      .A1(execution_unit_0_alu_0_n_49_1), .A2(execution_unit_0_alu_out[2]), .A3(
      execution_unit_0_alu_out[3]), .A4(execution_unit_0_alu_out[4]));
  OR3_X1_LVT execution_unit_0_alu_0_i_49_3 (.ZN(execution_unit_0_alu_0_n_49_3), 
      .A1(execution_unit_0_alu_0_n_49_2), .A2(execution_unit_0_alu_out[0]), .A3(
      execution_unit_0_alu_out[1]));
  NOR4_X1_LVT execution_unit_0_alu_0_i_49_4 (.ZN(execution_unit_0_alu_0_n_49_4), 
      .A1(execution_unit_0_alu_out[13]), .A2(execution_unit_0_alu_out[14]), .A3(
      execution_unit_0_alu_out[15]), .A4(inst_bw));
  NOR4_X1_LVT execution_unit_0_alu_0_i_49_5 (.ZN(execution_unit_0_alu_0_n_49_5), 
      .A1(execution_unit_0_alu_out[5]), .A2(execution_unit_0_alu_out[6]), .A3(
      execution_unit_0_alu_out[7]), .A4(execution_unit_0_alu_out[8]));
  NOR4_X1_LVT execution_unit_0_alu_0_i_49_6 (.ZN(execution_unit_0_alu_0_n_49_6), 
      .A1(execution_unit_0_alu_out[9]), .A2(execution_unit_0_alu_out[10]), .A3(
      execution_unit_0_alu_out[11]), .A4(execution_unit_0_alu_out[12]));
  INV_X1_LVT execution_unit_0_alu_0_i_49_7 (.ZN(execution_unit_0_alu_0_n_49_7), 
      .A(execution_unit_0_alu_out[4]));
  NAND4_X1_LVT execution_unit_0_alu_0_i_49_8 (.ZN(execution_unit_0_alu_0_n_49_8), 
      .A1(execution_unit_0_alu_0_n_49_4), .A2(execution_unit_0_alu_0_n_49_5), 
      .A3(execution_unit_0_alu_0_n_49_6), .A4(execution_unit_0_alu_0_n_49_7));
  OR4_X1_LVT execution_unit_0_alu_0_i_49_9 (.ZN(execution_unit_0_alu_0_n_49_9), 
      .A1(execution_unit_0_alu_0_n_49_8), .A2(execution_unit_0_alu_out[1]), .A3(
      execution_unit_0_alu_out[2]), .A4(execution_unit_0_alu_out[3]));
  OAI21_X1_LVT execution_unit_0_alu_0_i_49_10 (.ZN(execution_unit_0_alu_0_Z), .A(
      execution_unit_0_alu_0_n_49_3), .B1(execution_unit_0_alu_0_n_49_9), .B2(
      execution_unit_0_alu_out[0]));
  INV_X1_LVT execution_unit_0_alu_0_i_50_0 (.ZN(execution_unit_0_alu_0_n_112), 
      .A(execution_unit_0_alu_0_Z));
  NAND2_X1_LVT execution_unit_0_alu_0_i_51_5 (.ZN(execution_unit_0_alu_0_n_51_5), 
      .A1(execution_unit_0_alu_0_n_51_4), .A2(execution_unit_0_alu_0_n_112));
  XNOR2_X1_LVT execution_unit_0_alu_0_i_41_16 (.ZN(
      execution_unit_0_alu_0_n_41_16), .A(execution_unit_0_alu_0_alu_add[16]), 
      .B(execution_unit_0_alu_0_n_41_15));
  INV_X1_LVT execution_unit_0_alu_0_i_41_17 (.ZN(
      execution_unit_0_alu_0_alu_add_inc[16]), .A(execution_unit_0_alu_0_n_41_16));
  OR2_X1_LVT execution_unit_0_alu_0_i_27_7 (.ZN(execution_unit_0_alu_0_n_27_5), 
      .A1(execution_unit_0_alu_0_n_82), .A2(execution_unit_0_alu_0_n_84));
  HA_X1_LVT execution_unit_0_alu_0_i_26_2 (.CO(execution_unit_0_alu_0_n_26_2), 
      .S(execution_unit_0_alu_0_n_85), .A(execution_unit_0_alu_0_n_80), .B(
      execution_unit_0_alu_0_n_26_1));
  INV_X1_LVT execution_unit_0_alu_0_i_27_8 (.ZN(execution_unit_0_alu_0_n_27_6), 
      .A(execution_unit_0_alu_0_n_85));
  XNOR2_X1_LVT execution_unit_0_alu_0_i_27_10 (.ZN(execution_unit_0_alu_0_n_27_8), 
      .A(execution_unit_0_alu_0_n_27_5), .B(execution_unit_0_alu_0_n_27_6));
  XNOR2_X1_LVT execution_unit_0_alu_0_i_27_11 (.ZN(
      execution_unit_0_alu_0_bcd_add2[4]), .A(execution_unit_0_alu_0_n_27_8), .B(
      execution_unit_0_alu_0_n_27_7));
  AOI22_X1_LVT execution_unit_0_alu_0_i_44_32 (.ZN(
      execution_unit_0_alu_0_n_44_16), .A1(execution_unit_0_alu_0_n_104), .A2(
      execution_unit_0_alu_0_alu_add_inc[16]), .B1(execution_unit_0_alu_0_n_106), 
      .B2(execution_unit_0_alu_0_bcd_add2[4]));
  INV_X1_LVT execution_unit_0_alu_0_i_44_33 (.ZN(execution_unit_0_alu_0_n_107), 
      .A(execution_unit_0_alu_0_n_44_16));
  AOI22_X1_LVT execution_unit_0_alu_0_i_51_9 (.ZN(execution_unit_0_alu_0_n_51_9), 
      .A1(execution_unit_0_alu_0_n_51_8), .A2(execution_unit_0_alu_0_n_107), .B1(
      execution_unit_0_alu_out[8]), .B2(inst_bw));
  OAI211_X1_LVT execution_unit_0_alu_0_i_51_10 (.ZN(execution_unit_0_alu_stat[0]), 
      .A(execution_unit_0_alu_0_n_51_0), .B(execution_unit_0_alu_0_n_51_5), .C1(
      execution_unit_0_alu_0_n_51_7), .C2(execution_unit_0_alu_0_n_51_9));
  AND2_X1_LVT execution_unit_0_alu_0_i_52_0 (.ZN(execution_unit_0_alu_stat_wr[0]), 
      .A1(inst_alu[9]), .A2(execution_unit_0_n_0));
  NAND3_X1_LVT execution_unit_0_i_21_0 (.ZN(execution_unit_0_n_21_0), .A1(
      inst_type[2]), .A2(inst_ad[0]), .A3(execution_unit_0_n_13));
  NAND3_X1_LVT execution_unit_0_i_21_1 (.ZN(execution_unit_0_n_21_1), .A1(
      inst_as[0]), .A2(execution_unit_0_n_39), .A3(inst_type[0]));
  INV_X1_LVT execution_unit_0_i_21_2 (.ZN(execution_unit_0_n_21_2), .A(
      inst_type[1]));
  NAND3_X1_LVT execution_unit_0_i_21_3 (.ZN(execution_unit_0_n_21_3), .A1(
      execution_unit_0_n_21_0), .A2(execution_unit_0_n_21_1), .A3(
      execution_unit_0_n_21_2));
  AOI21_X1_LVT execution_unit_0_i_21_4 (.ZN(execution_unit_0_n_21_4), .A(
      dbg_reg_wr), .B1(execution_unit_0_n_21_3), .B2(execution_unit_0_n_0));
  INV_X1_LVT execution_unit_0_i_21_5 (.ZN(execution_unit_0_reg_dest_wr), .A(
      execution_unit_0_n_21_4));
  AOI21_X1_LVT execution_unit_0_i_23_0 (.ZN(execution_unit_0_n_23_0), .A(
      execution_unit_0_n_40), .B1(inst_so[5]), .B2(execution_unit_0_n_0));
  INV_X1_LVT execution_unit_0_i_23_1 (.ZN(execution_unit_0_reg_pc_call), .A(
      execution_unit_0_n_23_0));
  AND2_X1_LVT execution_unit_0_i_30_0 (.ZN(execution_unit_0_n_30_0), .A1(
      execution_unit_0_n_11), .A2(execution_unit_0_n_46));
  INV_X1_LVT execution_unit_0_i_30_1 (.ZN(execution_unit_0_n_30_1), .A(
      execution_unit_0_n_45));
  NOR3_X1_LVT execution_unit_0_i_30_2 (.ZN(execution_unit_0_n_30_2), .A1(
      execution_unit_0_n_30_1), .A2(execution_unit_0_n_42), .A3(inst_as[1]));
  OR4_X1_LVT execution_unit_0_i_30_3 (.ZN(execution_unit_0_reg_sp_wr), .A1(
      execution_unit_0_n_30_0), .A2(execution_unit_0_n_30_2), .A3(
      execution_unit_0_n_44), .A4(execution_unit_0_n_43));
  AOI221_X1_LVT execution_unit_0_i_32_0 (.ZN(execution_unit_0_n_32_0), .A(
      execution_unit_0_n_9), .B1(exec_done), .B2(inst_as[3]), .C1(
      execution_unit_0_n_1), .C2(inst_so[6]));
  INV_X1_LVT execution_unit_0_i_32_1 (.ZN(execution_unit_0_reg_incr), .A(
      execution_unit_0_n_32_0));
  INV_X1_LVT execution_unit_0_register_file_0_i_6_0 (.ZN(
      execution_unit_0_register_file_0_n_6_0), .A(execution_unit_0_reg_sr_clr));
  AOI21_X1_LVT execution_unit_0_register_file_0_i_1_0 (.ZN(
      execution_unit_0_register_file_0_n_1_0), .A(execution_unit_0_reg_sr_wr), 
      .B1(inst_dest[2]), .B2(execution_unit_0_reg_dest_wr));
  INV_X1_LVT execution_unit_0_register_file_0_i_1_1 (.ZN(
      execution_unit_0_register_file_0_r2_wr), .A(
      execution_unit_0_register_file_0_n_1_0));
  INV_X1_LVT execution_unit_0_register_file_0_i_2_0 (.ZN(
      execution_unit_0_register_file_0_n_2_0), .A(
      execution_unit_0_register_file_0_r2_wr));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_2_3 (.ZN(
      execution_unit_0_register_file_0_n_2_2), .A1(
      execution_unit_0_register_file_0_n_2_0), .A2(
      execution_unit_0_register_file_0_n_7), .B1(
      execution_unit_0_register_file_0_r2_wr), .B2(execution_unit_0_alu_out[4]));
  INV_X1_LVT execution_unit_0_register_file_0_i_2_4 (.ZN(
      execution_unit_0_register_file_0_r2_nxt[1]), .A(
      execution_unit_0_register_file_0_n_2_2));
  AND2_X1_LVT execution_unit_0_register_file_0_i_6_5 (.ZN(
      execution_unit_0_register_file_0_n_17), .A1(
      execution_unit_0_register_file_0_n_6_0), .A2(
      execution_unit_0_register_file_0_r2_nxt[1]));
  INV_X1_LVT execution_unit_0_register_file_0_i_3_0 (.ZN(
      execution_unit_0_register_file_0_n_8), .A(puc_rst));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r2_reg[4] (.Q(
      execution_unit_0_register_file_0_n_7), .QN(), .CK(cpu_mclk), .D(
      execution_unit_0_register_file_0_n_17), .RN(
      execution_unit_0_register_file_0_n_8));
  AOI21_X1_LVT execution_unit_0_register_file_0_i_8_0 (.ZN(
      execution_unit_0_register_file_0_n_8_0), .A(
      execution_unit_0_register_file_0_n_7), .B1(
      execution_unit_0_register_file_0_r2_nxt[1]), .B2(
      execution_unit_0_register_file_0_r2_wr));
  INV_X1_LVT execution_unit_0_register_file_0_i_8_1 (.ZN(cpuoff), .A(
      execution_unit_0_register_file_0_n_8_0));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_2_1 (.ZN(
      execution_unit_0_register_file_0_n_2_1), .A1(
      execution_unit_0_register_file_0_n_2_0), .A2(gie), .B1(
      execution_unit_0_alu_out[3]), .B2(execution_unit_0_register_file_0_r2_wr));
  INV_X1_LVT execution_unit_0_register_file_0_i_2_2 (.ZN(
      execution_unit_0_register_file_0_r2_nxt[0]), .A(
      execution_unit_0_register_file_0_n_2_1));
  AND2_X1_LVT execution_unit_0_register_file_0_i_6_4 (.ZN(
      execution_unit_0_register_file_0_n_16), .A1(
      execution_unit_0_register_file_0_n_6_0), .A2(
      execution_unit_0_register_file_0_r2_nxt[0]));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r2_reg[3] (.Q(gie), .QN(), .CK(
      cpu_mclk), .D(execution_unit_0_register_file_0_n_16), .RN(
      execution_unit_0_register_file_0_n_8));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r2_reg[5] (.Q(oscoff), .QN(), 
      .CK(cpu_mclk), .D(1'b0), .RN(execution_unit_0_register_file_0_n_8));
  INV_X1_LVT execution_unit_0_register_file_0_i_0_0 (.ZN(
      execution_unit_0_register_file_0_n_0_0), .A(inst_bw));
  AND2_X1_LVT execution_unit_0_register_file_0_i_0_8 (.ZN(pc_sw[15]), .A1(
      execution_unit_0_register_file_0_n_0_0), .A2(execution_unit_0_alu_out[15]));
  AND2_X1_LVT execution_unit_0_register_file_0_i_0_7 (.ZN(pc_sw[14]), .A1(
      execution_unit_0_register_file_0_n_0_0), .A2(execution_unit_0_alu_out[14]));
  AND2_X1_LVT execution_unit_0_register_file_0_i_0_6 (.ZN(pc_sw[13]), .A1(
      execution_unit_0_register_file_0_n_0_0), .A2(execution_unit_0_alu_out[13]));
  AND2_X1_LVT execution_unit_0_register_file_0_i_0_5 (.ZN(pc_sw[12]), .A1(
      execution_unit_0_register_file_0_n_0_0), .A2(execution_unit_0_alu_out[12]));
  AND2_X1_LVT execution_unit_0_register_file_0_i_0_4 (.ZN(pc_sw[11]), .A1(
      execution_unit_0_register_file_0_n_0_0), .A2(execution_unit_0_alu_out[11]));
  AND2_X1_LVT execution_unit_0_register_file_0_i_0_3 (.ZN(pc_sw[10]), .A1(
      execution_unit_0_register_file_0_n_0_0), .A2(execution_unit_0_alu_out[10]));
  AND2_X1_LVT execution_unit_0_register_file_0_i_0_2 (.ZN(pc_sw[9]), .A1(
      execution_unit_0_register_file_0_n_0_0), .A2(execution_unit_0_alu_out[9]));
  AND2_X1_LVT execution_unit_0_register_file_0_i_0_1 (.ZN(pc_sw[8]), .A1(
      execution_unit_0_register_file_0_n_0_0), .A2(execution_unit_0_alu_out[8]));
  AOI21_X1_LVT execution_unit_0_register_file_0_i_9_0 (.ZN(
      execution_unit_0_register_file_0_n_9_0), .A(execution_unit_0_reg_pc_call), 
      .B1(inst_dest[0]), .B2(execution_unit_0_reg_dest_wr));
  INV_X1_LVT execution_unit_0_register_file_0_i_9_1 (.ZN(pc_sw_wr), .A(
      execution_unit_0_register_file_0_n_9_0));
  AND2_X1_LVT execution_unit_0_register_file_0_i_19_0 (.ZN(
      execution_unit_0_register_file_0_r4_wr), .A1(inst_dest[4]), .A2(
      execution_unit_0_reg_dest_wr));
  INV_X1_LVT execution_unit_0_register_file_0_i_24_0 (.ZN(
      execution_unit_0_register_file_0_n_24_0), .A(
      execution_unit_0_register_file_0_r4_wr));
  INV_X1_LVT execution_unit_0_register_file_0_i_17_0 (.ZN(
      execution_unit_0_register_file_0_n_17_0), .A(inst_src[4]));
  NOR2_X1_LVT execution_unit_0_register_file_0_i_17_1 (.ZN(
      execution_unit_0_register_file_0_n_24), .A1(
      execution_unit_0_register_file_0_n_17_0), .A2(execution_unit_0_reg_sr_clr));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_315 (.ZN(
      execution_unit_0_register_file_0_n_105_300), .A1(
      execution_unit_0_register_file_0_n_24), .A2(
      execution_unit_0_register_file_0_r4[15]));
  INV_X1_LVT execution_unit_0_register_file_0_i_14_0 (.ZN(
      execution_unit_0_register_file_0_n_14_0), .A(inst_src[3]));
  NOR2_X1_LVT execution_unit_0_register_file_0_i_14_1 (.ZN(
      execution_unit_0_register_file_0_n_22), .A1(
      execution_unit_0_register_file_0_n_14_0), .A2(execution_unit_0_reg_sr_clr));
  AND2_X1_LVT execution_unit_0_register_file_0_i_15_0 (.ZN(
      execution_unit_0_register_file_0_r3_wr), .A1(inst_dest[3]), .A2(
      execution_unit_0_reg_dest_wr));
  CLKGATETST_X1_LVT execution_unit_0_register_file_0_clk_gate_r3_reg (.GCK(
      execution_unit_0_register_file_0_n_23), .CK(cpu_mclk), .E(
      execution_unit_0_register_file_0_r3_wr), .SE(1'b0));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r3_reg[15] (.Q(
      execution_unit_0_register_file_0_r3[15]), .QN(), .CK(
      execution_unit_0_register_file_0_n_23), .D(pc_sw[15]), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_316 (.ZN(
      execution_unit_0_register_file_0_n_105_301), .A1(
      execution_unit_0_register_file_0_n_22), .A2(
      execution_unit_0_register_file_0_r3[15]));
  INV_X1_LVT execution_unit_0_register_file_0_i_13_1 (.ZN(
      execution_unit_0_register_file_0_n_13_1), .A(inst_src[2]));
  INV_X1_LVT execution_unit_0_register_file_0_i_13_0 (.ZN(
      execution_unit_0_register_file_0_n_13_0), .A(execution_unit_0_reg_sr_clr));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_13_2 (.ZN(
      execution_unit_0_register_file_0_n_21), .A1(
      execution_unit_0_register_file_0_n_13_1), .A2(
      execution_unit_0_register_file_0_n_13_0));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r2_reg[15] (.Q(
      execution_unit_0_register_file_0_n_0), .QN(), .CK(cpu_mclk), .D(1'b0), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_317 (.ZN(
      execution_unit_0_register_file_0_n_105_302), .A1(
      execution_unit_0_register_file_0_n_21), .A2(
      execution_unit_0_register_file_0_n_0));
  INV_X1_LVT execution_unit_0_register_file_0_i_10_0 (.ZN(
      execution_unit_0_register_file_0_n_10_0), .A(inst_src[1]));
  NOR2_X1_LVT execution_unit_0_register_file_0_i_10_1 (.ZN(
      execution_unit_0_register_file_0_inst_src_in), .A1(
      execution_unit_0_register_file_0_n_10_0), .A2(execution_unit_0_reg_sr_clr));
  AND2_X1_LVT execution_unit_0_register_file_0_i_12_0 (.ZN(
      execution_unit_0_register_file_0_r1_wr), .A1(inst_dest[1]), .A2(
      execution_unit_0_reg_dest_wr));
  INV_X1_LVT execution_unit_0_register_file_0_i_108_1 (.ZN(
      execution_unit_0_register_file_0_n_108_0), .A(execution_unit_0_reg_sp_wr));
  NOR2_X1_LVT execution_unit_0_register_file_0_i_108_2 (.ZN(
      execution_unit_0_register_file_0_n_272), .A1(
      execution_unit_0_register_file_0_n_108_0), .A2(
      execution_unit_0_register_file_0_r1_wr));
  NOR2_X1_LVT execution_unit_0_register_file_0_i_108_0 (.ZN(
      execution_unit_0_register_file_0_n_271), .A1(execution_unit_0_reg_sp_wr), 
      .A2(execution_unit_0_register_file_0_r1_wr));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_24_27 (.ZN(
      execution_unit_0_register_file_0_n_24_14), .A1(
      execution_unit_0_register_file_0_n_24_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[13]), .B1(
      execution_unit_0_register_file_0_r4_wr), .B2(pc_sw[13]));
  INV_X1_LVT execution_unit_0_register_file_0_i_24_28 (.ZN(
      execution_unit_0_register_file_0_n_41), .A(
      execution_unit_0_register_file_0_n_24_14));
  AND2_X1_LVT execution_unit_0_register_file_0_i_18_0 (.ZN(
      execution_unit_0_register_file_0_r4_inc), .A1(
      execution_unit_0_register_file_0_n_24), .A2(execution_unit_0_reg_incr));
  INV_X1_LVT execution_unit_0_register_file_0_i_25_1 (.ZN(
      execution_unit_0_register_file_0_n_25_1), .A(
      execution_unit_0_register_file_0_r4_inc));
  INV_X1_LVT execution_unit_0_register_file_0_i_25_0 (.ZN(
      execution_unit_0_register_file_0_n_25_0), .A(
      execution_unit_0_register_file_0_r4_wr));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_25_2 (.ZN(
      execution_unit_0_register_file_0_n_44), .A1(
      execution_unit_0_register_file_0_n_25_1), .A2(
      execution_unit_0_register_file_0_n_25_0));
  CLKGATETST_X1_LVT execution_unit_0_register_file_0_clk_gate_r4_reg (.GCK(
      execution_unit_0_register_file_0_n_27), .CK(cpu_mclk), .E(
      execution_unit_0_register_file_0_n_44), .SE(1'b0));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r4_reg[13] (.Q(
      execution_unit_0_register_file_0_r4[13]), .QN(), .CK(
      execution_unit_0_register_file_0_n_27), .D(
      execution_unit_0_register_file_0_n_41), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_273 (.ZN(
      execution_unit_0_register_file_0_n_105_260), .A1(
      execution_unit_0_register_file_0_n_24), .A2(
      execution_unit_0_register_file_0_r4[13]));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r3_reg[13] (.Q(
      execution_unit_0_register_file_0_r3[13]), .QN(), .CK(
      execution_unit_0_register_file_0_n_23), .D(pc_sw[13]), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_274 (.ZN(
      execution_unit_0_register_file_0_n_105_261), .A1(
      execution_unit_0_register_file_0_n_22), .A2(
      execution_unit_0_register_file_0_r3[13]));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r2_reg[13] (.Q(
      execution_unit_0_register_file_0_n_2), .QN(), .CK(cpu_mclk), .D(1'b0), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_275 (.ZN(
      execution_unit_0_register_file_0_n_105_262), .A1(
      execution_unit_0_register_file_0_n_21), .A2(
      execution_unit_0_register_file_0_n_2));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_24_23 (.ZN(
      execution_unit_0_register_file_0_n_24_12), .A1(
      execution_unit_0_register_file_0_n_24_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[11]), .B1(
      execution_unit_0_register_file_0_r4_wr), .B2(pc_sw[11]));
  INV_X1_LVT execution_unit_0_register_file_0_i_24_24 (.ZN(
      execution_unit_0_register_file_0_n_39), .A(
      execution_unit_0_register_file_0_n_24_12));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r4_reg[11] (.Q(
      execution_unit_0_register_file_0_r4[11]), .QN(), .CK(
      execution_unit_0_register_file_0_n_27), .D(
      execution_unit_0_register_file_0_n_39), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_231 (.ZN(
      execution_unit_0_register_file_0_n_105_220), .A1(
      execution_unit_0_register_file_0_n_24), .A2(
      execution_unit_0_register_file_0_r4[11]));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r3_reg[11] (.Q(
      execution_unit_0_register_file_0_r3[11]), .QN(), .CK(
      execution_unit_0_register_file_0_n_23), .D(pc_sw[11]), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_232 (.ZN(
      execution_unit_0_register_file_0_n_105_221), .A1(
      execution_unit_0_register_file_0_n_22), .A2(
      execution_unit_0_register_file_0_r3[11]));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r2_reg[11] (.Q(
      execution_unit_0_register_file_0_n_4), .QN(), .CK(cpu_mclk), .D(1'b0), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_233 (.ZN(
      execution_unit_0_register_file_0_n_105_222), .A1(
      execution_unit_0_register_file_0_n_21), .A2(
      execution_unit_0_register_file_0_n_4));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_24_19 (.ZN(
      execution_unit_0_register_file_0_n_24_10), .A1(
      execution_unit_0_register_file_0_n_24_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[9]), .B1(
      execution_unit_0_register_file_0_r4_wr), .B2(pc_sw[9]));
  INV_X1_LVT execution_unit_0_register_file_0_i_24_20 (.ZN(
      execution_unit_0_register_file_0_n_37), .A(
      execution_unit_0_register_file_0_n_24_10));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r4_reg[9] (.Q(
      execution_unit_0_register_file_0_r4[9]), .QN(), .CK(
      execution_unit_0_register_file_0_n_27), .D(
      execution_unit_0_register_file_0_n_37), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_189 (.ZN(
      execution_unit_0_register_file_0_n_105_180), .A1(
      execution_unit_0_register_file_0_n_24), .A2(
      execution_unit_0_register_file_0_r4[9]));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r3_reg[9] (.Q(
      execution_unit_0_register_file_0_r3[9]), .QN(), .CK(
      execution_unit_0_register_file_0_n_23), .D(pc_sw[9]), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_190 (.ZN(
      execution_unit_0_register_file_0_n_105_181), .A1(
      execution_unit_0_register_file_0_n_22), .A2(
      execution_unit_0_register_file_0_r3[9]));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r2_reg[9] (.Q(
      execution_unit_0_register_file_0_n_6), .QN(), .CK(cpu_mclk), .D(1'b0), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_191 (.ZN(
      execution_unit_0_register_file_0_n_105_182), .A1(
      execution_unit_0_register_file_0_n_21), .A2(
      execution_unit_0_register_file_0_n_6));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_24_15 (.ZN(
      execution_unit_0_register_file_0_n_24_8), .A1(
      execution_unit_0_register_file_0_n_24_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[7]), .B1(
      execution_unit_0_register_file_0_r4_wr), .B2(execution_unit_0_alu_out[7]));
  INV_X1_LVT execution_unit_0_register_file_0_i_24_16 (.ZN(
      execution_unit_0_register_file_0_n_35), .A(
      execution_unit_0_register_file_0_n_24_8));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r4_reg[7] (.Q(
      execution_unit_0_register_file_0_r4[7]), .QN(), .CK(
      execution_unit_0_register_file_0_n_27), .D(
      execution_unit_0_register_file_0_n_35), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_147 (.ZN(
      execution_unit_0_register_file_0_n_105_140), .A1(
      execution_unit_0_register_file_0_n_24), .A2(
      execution_unit_0_register_file_0_r4[7]));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r3_reg[7] (.Q(
      execution_unit_0_register_file_0_r3[7]), .QN(), .CK(
      execution_unit_0_register_file_0_n_23), .D(execution_unit_0_alu_out[7]), 
      .RN(execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_148 (.ZN(
      execution_unit_0_register_file_0_n_105_141), .A1(
      execution_unit_0_register_file_0_n_22), .A2(
      execution_unit_0_register_file_0_r3[7]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_2_7 (.ZN(
      execution_unit_0_register_file_0_n_2_4), .A1(
      execution_unit_0_register_file_0_n_2_0), .A2(scg1), .B1(
      execution_unit_0_register_file_0_r2_wr), .B2(execution_unit_0_alu_out[7]));
  INV_X1_LVT execution_unit_0_register_file_0_i_2_8 (.ZN(
      execution_unit_0_register_file_0_r2_nxt[4]), .A(
      execution_unit_0_register_file_0_n_2_4));
  AND2_X1_LVT execution_unit_0_register_file_0_i_6_7 (.ZN(
      execution_unit_0_register_file_0_n_19), .A1(
      execution_unit_0_register_file_0_n_6_0), .A2(
      execution_unit_0_register_file_0_r2_nxt[4]));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r2_reg[7] (.Q(scg1), .QN(), .CK(
      cpu_mclk), .D(execution_unit_0_register_file_0_n_19), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_149 (.ZN(
      execution_unit_0_register_file_0_n_105_142), .A1(
      execution_unit_0_register_file_0_n_21), .A2(scg1));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_24_11 (.ZN(
      execution_unit_0_register_file_0_n_24_6), .A1(
      execution_unit_0_register_file_0_n_24_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[5]), .B1(
      execution_unit_0_register_file_0_r4_wr), .B2(execution_unit_0_alu_out[5]));
  INV_X1_LVT execution_unit_0_register_file_0_i_24_12 (.ZN(
      execution_unit_0_register_file_0_n_33), .A(
      execution_unit_0_register_file_0_n_24_6));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r4_reg[5] (.Q(
      execution_unit_0_register_file_0_r4[5]), .QN(), .CK(
      execution_unit_0_register_file_0_n_27), .D(
      execution_unit_0_register_file_0_n_33), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_105 (.ZN(
      execution_unit_0_register_file_0_n_105_100), .A1(
      execution_unit_0_register_file_0_n_24), .A2(
      execution_unit_0_register_file_0_r4[5]));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r3_reg[5] (.Q(
      execution_unit_0_register_file_0_r3[5]), .QN(), .CK(
      execution_unit_0_register_file_0_n_23), .D(execution_unit_0_alu_out[5]), 
      .RN(execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_106 (.ZN(
      execution_unit_0_register_file_0_n_105_101), .A1(
      execution_unit_0_register_file_0_n_22), .A2(
      execution_unit_0_register_file_0_r3[5]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_107 (.ZN(
      execution_unit_0_register_file_0_n_105_102), .A1(
      execution_unit_0_register_file_0_n_21), .A2(oscoff));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_24_7 (.ZN(
      execution_unit_0_register_file_0_n_24_4), .A1(
      execution_unit_0_register_file_0_n_24_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[3]), .B1(
      execution_unit_0_register_file_0_r4_wr), .B2(execution_unit_0_alu_out[3]));
  INV_X1_LVT execution_unit_0_register_file_0_i_24_8 (.ZN(
      execution_unit_0_register_file_0_n_31), .A(
      execution_unit_0_register_file_0_n_24_4));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r4_reg[3] (.Q(
      execution_unit_0_register_file_0_r4[3]), .QN(), .CK(
      execution_unit_0_register_file_0_n_27), .D(
      execution_unit_0_register_file_0_n_31), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_63 (.ZN(
      execution_unit_0_register_file_0_n_105_60), .A1(
      execution_unit_0_register_file_0_n_24), .A2(
      execution_unit_0_register_file_0_r4[3]));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r3_reg[3] (.Q(
      execution_unit_0_register_file_0_r3[3]), .QN(), .CK(
      execution_unit_0_register_file_0_n_23), .D(execution_unit_0_alu_out[3]), 
      .RN(execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_64 (.ZN(
      execution_unit_0_register_file_0_n_105_61), .A1(
      execution_unit_0_register_file_0_n_22), .A2(
      execution_unit_0_register_file_0_r3[3]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_65 (.ZN(
      execution_unit_0_register_file_0_n_105_62), .A1(
      execution_unit_0_register_file_0_n_21), .A2(gie));
  INV_X1_LVT execution_unit_0_register_file_0_i_20_0 (.ZN(
      execution_unit_0_register_file_0_n_20_0), .A(inst_bw));
  NOR2_X1_LVT execution_unit_0_register_file_0_i_20_1 (.ZN(
      execution_unit_0_register_file_0_n_25), .A1(
      execution_unit_0_register_file_0_n_20_0), .A2(
      execution_unit_0_register_file_0_inst_src_in));
  INV_X1_LVT execution_unit_0_register_file_0_i_21_0 (.ZN(
      execution_unit_0_register_file_0_n_26), .A(
      execution_unit_0_register_file_0_n_25));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_24_3 (.ZN(
      execution_unit_0_register_file_0_n_24_2), .A1(
      execution_unit_0_register_file_0_n_24_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[1]), .B1(
      execution_unit_0_register_file_0_r4_wr), .B2(execution_unit_0_alu_out[1]));
  INV_X1_LVT execution_unit_0_register_file_0_i_24_4 (.ZN(
      execution_unit_0_register_file_0_n_29), .A(
      execution_unit_0_register_file_0_n_24_2));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r4_reg[1] (.Q(
      execution_unit_0_register_file_0_r4[1]), .QN(), .CK(
      execution_unit_0_register_file_0_n_27), .D(
      execution_unit_0_register_file_0_n_29), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_21 (.ZN(
      execution_unit_0_register_file_0_n_105_20), .A1(
      execution_unit_0_register_file_0_n_24), .A2(
      execution_unit_0_register_file_0_r4[1]));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r3_reg[1] (.Q(
      execution_unit_0_register_file_0_r3[1]), .QN(), .CK(
      execution_unit_0_register_file_0_n_23), .D(execution_unit_0_alu_out[1]), 
      .RN(execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_22 (.ZN(
      execution_unit_0_register_file_0_n_105_21), .A1(
      execution_unit_0_register_file_0_n_22), .A2(
      execution_unit_0_register_file_0_r3[1]));
  INV_X1_LVT execution_unit_0_register_file_0_i_5_0 (.ZN(
      execution_unit_0_register_file_0_n_5_0), .A(
      execution_unit_0_register_file_0_r2_wr));
  INV_X1_LVT execution_unit_0_register_file_0_i_5_6 (.ZN(
      execution_unit_0_register_file_0_n_5_5), .A(
      execution_unit_0_alu_stat_wr[1]));
  NAND3_X1_LVT execution_unit_0_register_file_0_i_5_7 (.ZN(
      execution_unit_0_register_file_0_n_5_6), .A1(
      execution_unit_0_register_file_0_n_5_0), .A2(
      execution_unit_0_register_file_0_n_5_5), .A3(execution_unit_0_status[1]));
  NAND3_X1_LVT execution_unit_0_register_file_0_i_5_8 (.ZN(
      execution_unit_0_register_file_0_n_5_7), .A1(
      execution_unit_0_register_file_0_n_5_5), .A2(
      execution_unit_0_register_file_0_r2_wr), .A3(execution_unit_0_alu_out[1]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_5_9 (.ZN(
      execution_unit_0_register_file_0_n_5_8), .A1(execution_unit_0_alu_stat[1]), 
      .A2(execution_unit_0_alu_stat_wr[1]));
  NAND3_X1_LVT execution_unit_0_register_file_0_i_5_10 (.ZN(
      execution_unit_0_register_file_0_n_10), .A1(
      execution_unit_0_register_file_0_n_5_6), .A2(
      execution_unit_0_register_file_0_n_5_7), .A3(
      execution_unit_0_register_file_0_n_5_8));
  AND2_X1_LVT execution_unit_0_register_file_0_i_6_2 (.ZN(
      execution_unit_0_register_file_0_n_14), .A1(
      execution_unit_0_register_file_0_n_6_0), .A2(
      execution_unit_0_register_file_0_n_10));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r2_reg[1] (.Q(
      execution_unit_0_status[1]), .QN(), .CK(cpu_mclk), .D(
      execution_unit_0_register_file_0_n_14), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_23 (.ZN(
      execution_unit_0_register_file_0_n_105_22), .A1(
      execution_unit_0_register_file_0_n_21), .A2(execution_unit_0_status[1]));
  INV_X1_LVT execution_unit_0_register_file_0_i_106_0 (.ZN(
      execution_unit_0_register_file_0_n_255), .A(execution_unit_0_reg_src[1]));
  AOI222_X1_LVT execution_unit_0_register_file_0_i_109_0 (.ZN(
      execution_unit_0_register_file_0_n_109_0), .A1(
      execution_unit_0_register_file_0_r1_wr), .A2(execution_unit_0_alu_out[1]), 
      .B1(execution_unit_0_register_file_0_n_272), .B2(eu_mab[1]), .C1(
      execution_unit_0_register_file_0_n_271), .C2(
      execution_unit_0_register_file_0_n_255));
  INV_X1_LVT execution_unit_0_register_file_0_i_109_1 (.ZN(
      execution_unit_0_register_file_0_n_273), .A(
      execution_unit_0_register_file_0_n_109_0));
  INV_X1_LVT execution_unit_0_register_file_0_i_110_0 (.ZN(
      execution_unit_0_register_file_0_n_110_0), .A(execution_unit_0_reg_sp_wr));
  INV_X1_LVT execution_unit_0_register_file_0_i_110_1 (.ZN(
      execution_unit_0_register_file_0_n_110_1), .A(
      execution_unit_0_register_file_0_r1_wr));
  AND2_X1_LVT execution_unit_0_register_file_0_i_11_0 (.ZN(
      execution_unit_0_register_file_0_r1_inc), .A1(
      execution_unit_0_register_file_0_inst_src_in), .A2(
      execution_unit_0_reg_incr));
  NAND3_X1_LVT execution_unit_0_register_file_0_i_110_2 (.ZN(
      execution_unit_0_register_file_0_n_110_2), .A1(
      execution_unit_0_register_file_0_n_110_0), .A2(
      execution_unit_0_register_file_0_n_110_1), .A3(
      execution_unit_0_register_file_0_r1_inc));
  NAND3_X1_LVT execution_unit_0_register_file_0_i_110_3 (.ZN(
      execution_unit_0_register_file_0_n_288), .A1(
      execution_unit_0_register_file_0_n_110_2), .A2(
      execution_unit_0_register_file_0_n_110_0), .A3(
      execution_unit_0_register_file_0_n_110_1));
  CLKGATETST_X1_LVT execution_unit_0_register_file_0_clk_gate_r1_reg (.GCK(
      execution_unit_0_register_file_0_n_270), .CK(cpu_mclk), .E(
      execution_unit_0_register_file_0_n_288), .SE(1'b0));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r1_reg[1] (.Q(
      execution_unit_0_register_file_0_r1[1]), .QN(), .CK(
      execution_unit_0_register_file_0_n_270), .D(
      execution_unit_0_register_file_0_n_273), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_24 (.ZN(
      execution_unit_0_register_file_0_n_105_23), .A1(
      execution_unit_0_register_file_0_inst_src_in), .A2(
      execution_unit_0_register_file_0_r1[1]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_105_25 (.ZN(
      execution_unit_0_register_file_0_n_105_24), .A1(
      execution_unit_0_register_file_0_n_105_20), .A2(
      execution_unit_0_register_file_0_n_105_21), .A3(
      execution_unit_0_register_file_0_n_105_22), .A4(
      execution_unit_0_register_file_0_n_105_23));
  INV_X1_LVT execution_unit_0_register_file_0_i_76_0 (.ZN(
      execution_unit_0_register_file_0_n_76_0), .A(inst_src[12]));
  NOR2_X1_LVT execution_unit_0_register_file_0_i_76_1 (.ZN(
      execution_unit_0_register_file_0_n_178), .A1(
      execution_unit_0_register_file_0_n_76_0), .A2(execution_unit_0_reg_sr_clr));
  AND2_X1_LVT execution_unit_0_register_file_0_i_78_0 (.ZN(
      execution_unit_0_register_file_0_r12_wr), .A1(inst_dest[12]), .A2(
      execution_unit_0_reg_dest_wr));
  INV_X1_LVT execution_unit_0_register_file_0_i_80_0 (.ZN(
      execution_unit_0_register_file_0_n_80_0), .A(
      execution_unit_0_register_file_0_r12_wr));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_80_3 (.ZN(
      execution_unit_0_register_file_0_n_80_2), .A1(
      execution_unit_0_register_file_0_n_80_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[1]), .B1(
      execution_unit_0_register_file_0_r12_wr), .B2(execution_unit_0_alu_out[1]));
  INV_X1_LVT execution_unit_0_register_file_0_i_80_4 (.ZN(
      execution_unit_0_register_file_0_n_181), .A(
      execution_unit_0_register_file_0_n_80_2));
  AND2_X1_LVT execution_unit_0_register_file_0_i_77_0 (.ZN(
      execution_unit_0_register_file_0_r12_inc), .A1(
      execution_unit_0_register_file_0_n_178), .A2(execution_unit_0_reg_incr));
  INV_X1_LVT execution_unit_0_register_file_0_i_81_1 (.ZN(
      execution_unit_0_register_file_0_n_81_1), .A(
      execution_unit_0_register_file_0_r12_inc));
  INV_X1_LVT execution_unit_0_register_file_0_i_81_0 (.ZN(
      execution_unit_0_register_file_0_n_81_0), .A(
      execution_unit_0_register_file_0_r12_wr));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_81_2 (.ZN(
      execution_unit_0_register_file_0_n_196), .A1(
      execution_unit_0_register_file_0_n_81_1), .A2(
      execution_unit_0_register_file_0_n_81_0));
  CLKGATETST_X1_LVT execution_unit_0_register_file_0_clk_gate_r12_reg (.GCK(
      execution_unit_0_register_file_0_n_179), .CK(cpu_mclk), .E(
      execution_unit_0_register_file_0_n_196), .SE(1'b0));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r12_reg[1] (.Q(
      execution_unit_0_register_file_0_r12[1]), .QN(), .CK(
      execution_unit_0_register_file_0_n_179), .D(
      execution_unit_0_register_file_0_n_181), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_26 (.ZN(
      execution_unit_0_register_file_0_n_105_25), .A1(
      execution_unit_0_register_file_0_n_178), .A2(
      execution_unit_0_register_file_0_r12[1]));
  INV_X1_LVT execution_unit_0_register_file_0_i_69_0 (.ZN(
      execution_unit_0_register_file_0_n_69_0), .A(inst_src[11]));
  NOR2_X1_LVT execution_unit_0_register_file_0_i_69_1 (.ZN(
      execution_unit_0_register_file_0_n_159), .A1(
      execution_unit_0_register_file_0_n_69_0), .A2(execution_unit_0_reg_sr_clr));
  AND2_X1_LVT execution_unit_0_register_file_0_i_71_0 (.ZN(
      execution_unit_0_register_file_0_r11_wr), .A1(inst_dest[11]), .A2(
      execution_unit_0_reg_dest_wr));
  INV_X1_LVT execution_unit_0_register_file_0_i_73_0 (.ZN(
      execution_unit_0_register_file_0_n_73_0), .A(
      execution_unit_0_register_file_0_r11_wr));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_73_3 (.ZN(
      execution_unit_0_register_file_0_n_73_2), .A1(
      execution_unit_0_register_file_0_n_73_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[1]), .B1(
      execution_unit_0_register_file_0_r11_wr), .B2(execution_unit_0_alu_out[1]));
  INV_X1_LVT execution_unit_0_register_file_0_i_73_4 (.ZN(
      execution_unit_0_register_file_0_n_162), .A(
      execution_unit_0_register_file_0_n_73_2));
  AND2_X1_LVT execution_unit_0_register_file_0_i_70_0 (.ZN(
      execution_unit_0_register_file_0_r11_inc), .A1(
      execution_unit_0_register_file_0_n_159), .A2(execution_unit_0_reg_incr));
  INV_X1_LVT execution_unit_0_register_file_0_i_74_1 (.ZN(
      execution_unit_0_register_file_0_n_74_1), .A(
      execution_unit_0_register_file_0_r11_inc));
  INV_X1_LVT execution_unit_0_register_file_0_i_74_0 (.ZN(
      execution_unit_0_register_file_0_n_74_0), .A(
      execution_unit_0_register_file_0_r11_wr));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_74_2 (.ZN(
      execution_unit_0_register_file_0_n_177), .A1(
      execution_unit_0_register_file_0_n_74_1), .A2(
      execution_unit_0_register_file_0_n_74_0));
  CLKGATETST_X1_LVT execution_unit_0_register_file_0_clk_gate_r11_reg (.GCK(
      execution_unit_0_register_file_0_n_160), .CK(cpu_mclk), .E(
      execution_unit_0_register_file_0_n_177), .SE(1'b0));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r11_reg[1] (.Q(
      execution_unit_0_register_file_0_r11[1]), .QN(), .CK(
      execution_unit_0_register_file_0_n_160), .D(
      execution_unit_0_register_file_0_n_162), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_27 (.ZN(
      execution_unit_0_register_file_0_n_105_26), .A1(
      execution_unit_0_register_file_0_n_159), .A2(
      execution_unit_0_register_file_0_r11[1]));
  INV_X1_LVT execution_unit_0_register_file_0_i_62_0 (.ZN(
      execution_unit_0_register_file_0_n_62_0), .A(inst_src[10]));
  NOR2_X1_LVT execution_unit_0_register_file_0_i_62_1 (.ZN(
      execution_unit_0_register_file_0_n_140), .A1(
      execution_unit_0_register_file_0_n_62_0), .A2(execution_unit_0_reg_sr_clr));
  AND2_X1_LVT execution_unit_0_register_file_0_i_64_0 (.ZN(
      execution_unit_0_register_file_0_r10_wr), .A1(inst_dest[10]), .A2(
      execution_unit_0_reg_dest_wr));
  INV_X1_LVT execution_unit_0_register_file_0_i_66_0 (.ZN(
      execution_unit_0_register_file_0_n_66_0), .A(
      execution_unit_0_register_file_0_r10_wr));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_66_3 (.ZN(
      execution_unit_0_register_file_0_n_66_2), .A1(
      execution_unit_0_register_file_0_n_66_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[1]), .B1(
      execution_unit_0_register_file_0_r10_wr), .B2(execution_unit_0_alu_out[1]));
  INV_X1_LVT execution_unit_0_register_file_0_i_66_4 (.ZN(
      execution_unit_0_register_file_0_n_143), .A(
      execution_unit_0_register_file_0_n_66_2));
  AND2_X1_LVT execution_unit_0_register_file_0_i_63_0 (.ZN(
      execution_unit_0_register_file_0_r10_inc), .A1(
      execution_unit_0_register_file_0_n_140), .A2(execution_unit_0_reg_incr));
  INV_X1_LVT execution_unit_0_register_file_0_i_67_1 (.ZN(
      execution_unit_0_register_file_0_n_67_1), .A(
      execution_unit_0_register_file_0_r10_inc));
  INV_X1_LVT execution_unit_0_register_file_0_i_67_0 (.ZN(
      execution_unit_0_register_file_0_n_67_0), .A(
      execution_unit_0_register_file_0_r10_wr));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_67_2 (.ZN(
      execution_unit_0_register_file_0_n_158), .A1(
      execution_unit_0_register_file_0_n_67_1), .A2(
      execution_unit_0_register_file_0_n_67_0));
  CLKGATETST_X1_LVT execution_unit_0_register_file_0_clk_gate_r10_reg (.GCK(
      execution_unit_0_register_file_0_n_141), .CK(cpu_mclk), .E(
      execution_unit_0_register_file_0_n_158), .SE(1'b0));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r10_reg[1] (.Q(
      execution_unit_0_register_file_0_r10[1]), .QN(), .CK(
      execution_unit_0_register_file_0_n_141), .D(
      execution_unit_0_register_file_0_n_143), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_28 (.ZN(
      execution_unit_0_register_file_0_n_105_27), .A1(
      execution_unit_0_register_file_0_n_140), .A2(
      execution_unit_0_register_file_0_r10[1]));
  INV_X1_LVT execution_unit_0_register_file_0_i_55_0 (.ZN(
      execution_unit_0_register_file_0_n_55_0), .A(inst_src[9]));
  NOR2_X1_LVT execution_unit_0_register_file_0_i_55_1 (.ZN(
      execution_unit_0_register_file_0_n_121), .A1(
      execution_unit_0_register_file_0_n_55_0), .A2(execution_unit_0_reg_sr_clr));
  AND2_X1_LVT execution_unit_0_register_file_0_i_57_0 (.ZN(
      execution_unit_0_register_file_0_r9_wr), .A1(inst_dest[9]), .A2(
      execution_unit_0_reg_dest_wr));
  INV_X1_LVT execution_unit_0_register_file_0_i_59_0 (.ZN(
      execution_unit_0_register_file_0_n_59_0), .A(
      execution_unit_0_register_file_0_r9_wr));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_59_3 (.ZN(
      execution_unit_0_register_file_0_n_59_2), .A1(
      execution_unit_0_register_file_0_n_59_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[1]), .B1(
      execution_unit_0_register_file_0_r9_wr), .B2(execution_unit_0_alu_out[1]));
  INV_X1_LVT execution_unit_0_register_file_0_i_59_4 (.ZN(
      execution_unit_0_register_file_0_n_124), .A(
      execution_unit_0_register_file_0_n_59_2));
  AND2_X1_LVT execution_unit_0_register_file_0_i_56_0 (.ZN(
      execution_unit_0_register_file_0_r9_inc), .A1(
      execution_unit_0_register_file_0_n_121), .A2(execution_unit_0_reg_incr));
  INV_X1_LVT execution_unit_0_register_file_0_i_60_1 (.ZN(
      execution_unit_0_register_file_0_n_60_1), .A(
      execution_unit_0_register_file_0_r9_inc));
  INV_X1_LVT execution_unit_0_register_file_0_i_60_0 (.ZN(
      execution_unit_0_register_file_0_n_60_0), .A(
      execution_unit_0_register_file_0_r9_wr));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_60_2 (.ZN(
      execution_unit_0_register_file_0_n_139), .A1(
      execution_unit_0_register_file_0_n_60_1), .A2(
      execution_unit_0_register_file_0_n_60_0));
  CLKGATETST_X1_LVT execution_unit_0_register_file_0_clk_gate_r9_reg (.GCK(
      execution_unit_0_register_file_0_n_122), .CK(cpu_mclk), .E(
      execution_unit_0_register_file_0_n_139), .SE(1'b0));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r9_reg[1] (.Q(
      execution_unit_0_register_file_0_r9[1]), .QN(), .CK(
      execution_unit_0_register_file_0_n_122), .D(
      execution_unit_0_register_file_0_n_124), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_29 (.ZN(
      execution_unit_0_register_file_0_n_105_28), .A1(
      execution_unit_0_register_file_0_n_121), .A2(
      execution_unit_0_register_file_0_r9[1]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_105_30 (.ZN(
      execution_unit_0_register_file_0_n_105_29), .A1(
      execution_unit_0_register_file_0_n_105_25), .A2(
      execution_unit_0_register_file_0_n_105_26), .A3(
      execution_unit_0_register_file_0_n_105_27), .A4(
      execution_unit_0_register_file_0_n_105_28));
  INV_X1_LVT execution_unit_0_register_file_0_i_48_0 (.ZN(
      execution_unit_0_register_file_0_n_48_0), .A(inst_src[8]));
  NOR2_X1_LVT execution_unit_0_register_file_0_i_48_1 (.ZN(
      execution_unit_0_register_file_0_n_102), .A1(
      execution_unit_0_register_file_0_n_48_0), .A2(execution_unit_0_reg_sr_clr));
  AND2_X1_LVT execution_unit_0_register_file_0_i_50_0 (.ZN(
      execution_unit_0_register_file_0_r8_wr), .A1(inst_dest[8]), .A2(
      execution_unit_0_reg_dest_wr));
  INV_X1_LVT execution_unit_0_register_file_0_i_52_0 (.ZN(
      execution_unit_0_register_file_0_n_52_0), .A(
      execution_unit_0_register_file_0_r8_wr));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_52_3 (.ZN(
      execution_unit_0_register_file_0_n_52_2), .A1(
      execution_unit_0_register_file_0_n_52_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[1]), .B1(
      execution_unit_0_register_file_0_r8_wr), .B2(execution_unit_0_alu_out[1]));
  INV_X1_LVT execution_unit_0_register_file_0_i_52_4 (.ZN(
      execution_unit_0_register_file_0_n_105), .A(
      execution_unit_0_register_file_0_n_52_2));
  AND2_X1_LVT execution_unit_0_register_file_0_i_49_0 (.ZN(
      execution_unit_0_register_file_0_r8_inc), .A1(
      execution_unit_0_register_file_0_n_102), .A2(execution_unit_0_reg_incr));
  INV_X1_LVT execution_unit_0_register_file_0_i_53_1 (.ZN(
      execution_unit_0_register_file_0_n_53_1), .A(
      execution_unit_0_register_file_0_r8_inc));
  INV_X1_LVT execution_unit_0_register_file_0_i_53_0 (.ZN(
      execution_unit_0_register_file_0_n_53_0), .A(
      execution_unit_0_register_file_0_r8_wr));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_53_2 (.ZN(
      execution_unit_0_register_file_0_n_120), .A1(
      execution_unit_0_register_file_0_n_53_1), .A2(
      execution_unit_0_register_file_0_n_53_0));
  CLKGATETST_X1_LVT execution_unit_0_register_file_0_clk_gate_r8_reg (.GCK(
      execution_unit_0_register_file_0_n_103), .CK(cpu_mclk), .E(
      execution_unit_0_register_file_0_n_120), .SE(1'b0));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r8_reg[1] (.Q(
      execution_unit_0_register_file_0_r8[1]), .QN(), .CK(
      execution_unit_0_register_file_0_n_103), .D(
      execution_unit_0_register_file_0_n_105), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_31 (.ZN(
      execution_unit_0_register_file_0_n_105_30), .A1(
      execution_unit_0_register_file_0_n_102), .A2(
      execution_unit_0_register_file_0_r8[1]));
  INV_X1_LVT execution_unit_0_register_file_0_i_41_0 (.ZN(
      execution_unit_0_register_file_0_n_41_0), .A(inst_src[7]));
  NOR2_X1_LVT execution_unit_0_register_file_0_i_41_1 (.ZN(
      execution_unit_0_register_file_0_n_83), .A1(
      execution_unit_0_register_file_0_n_41_0), .A2(execution_unit_0_reg_sr_clr));
  AND2_X1_LVT execution_unit_0_register_file_0_i_43_0 (.ZN(
      execution_unit_0_register_file_0_r7_wr), .A1(inst_dest[7]), .A2(
      execution_unit_0_reg_dest_wr));
  INV_X1_LVT execution_unit_0_register_file_0_i_45_0 (.ZN(
      execution_unit_0_register_file_0_n_45_0), .A(
      execution_unit_0_register_file_0_r7_wr));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_45_3 (.ZN(
      execution_unit_0_register_file_0_n_45_2), .A1(
      execution_unit_0_register_file_0_n_45_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[1]), .B1(
      execution_unit_0_register_file_0_r7_wr), .B2(execution_unit_0_alu_out[1]));
  INV_X1_LVT execution_unit_0_register_file_0_i_45_4 (.ZN(
      execution_unit_0_register_file_0_n_86), .A(
      execution_unit_0_register_file_0_n_45_2));
  AND2_X1_LVT execution_unit_0_register_file_0_i_42_0 (.ZN(
      execution_unit_0_register_file_0_r7_inc), .A1(
      execution_unit_0_register_file_0_n_83), .A2(execution_unit_0_reg_incr));
  INV_X1_LVT execution_unit_0_register_file_0_i_46_1 (.ZN(
      execution_unit_0_register_file_0_n_46_1), .A(
      execution_unit_0_register_file_0_r7_inc));
  INV_X1_LVT execution_unit_0_register_file_0_i_46_0 (.ZN(
      execution_unit_0_register_file_0_n_46_0), .A(
      execution_unit_0_register_file_0_r7_wr));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_46_2 (.ZN(
      execution_unit_0_register_file_0_n_101), .A1(
      execution_unit_0_register_file_0_n_46_1), .A2(
      execution_unit_0_register_file_0_n_46_0));
  CLKGATETST_X1_LVT execution_unit_0_register_file_0_clk_gate_r7_reg (.GCK(
      execution_unit_0_register_file_0_n_84), .CK(cpu_mclk), .E(
      execution_unit_0_register_file_0_n_101), .SE(1'b0));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r7_reg[1] (.Q(
      execution_unit_0_register_file_0_r7[1]), .QN(), .CK(
      execution_unit_0_register_file_0_n_84), .D(
      execution_unit_0_register_file_0_n_86), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_32 (.ZN(
      execution_unit_0_register_file_0_n_105_31), .A1(
      execution_unit_0_register_file_0_n_83), .A2(
      execution_unit_0_register_file_0_r7[1]));
  INV_X1_LVT execution_unit_0_register_file_0_i_34_0 (.ZN(
      execution_unit_0_register_file_0_n_34_0), .A(inst_src[6]));
  NOR2_X1_LVT execution_unit_0_register_file_0_i_34_1 (.ZN(
      execution_unit_0_register_file_0_n_64), .A1(
      execution_unit_0_register_file_0_n_34_0), .A2(execution_unit_0_reg_sr_clr));
  AND2_X1_LVT execution_unit_0_register_file_0_i_36_0 (.ZN(
      execution_unit_0_register_file_0_r6_wr), .A1(inst_dest[6]), .A2(
      execution_unit_0_reg_dest_wr));
  INV_X1_LVT execution_unit_0_register_file_0_i_38_0 (.ZN(
      execution_unit_0_register_file_0_n_38_0), .A(
      execution_unit_0_register_file_0_r6_wr));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_38_3 (.ZN(
      execution_unit_0_register_file_0_n_38_2), .A1(
      execution_unit_0_register_file_0_n_38_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[1]), .B1(
      execution_unit_0_register_file_0_r6_wr), .B2(execution_unit_0_alu_out[1]));
  INV_X1_LVT execution_unit_0_register_file_0_i_38_4 (.ZN(
      execution_unit_0_register_file_0_n_67), .A(
      execution_unit_0_register_file_0_n_38_2));
  AND2_X1_LVT execution_unit_0_register_file_0_i_35_0 (.ZN(
      execution_unit_0_register_file_0_r6_inc), .A1(
      execution_unit_0_register_file_0_n_64), .A2(execution_unit_0_reg_incr));
  INV_X1_LVT execution_unit_0_register_file_0_i_39_1 (.ZN(
      execution_unit_0_register_file_0_n_39_1), .A(
      execution_unit_0_register_file_0_r6_inc));
  INV_X1_LVT execution_unit_0_register_file_0_i_39_0 (.ZN(
      execution_unit_0_register_file_0_n_39_0), .A(
      execution_unit_0_register_file_0_r6_wr));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_39_2 (.ZN(
      execution_unit_0_register_file_0_n_82), .A1(
      execution_unit_0_register_file_0_n_39_1), .A2(
      execution_unit_0_register_file_0_n_39_0));
  CLKGATETST_X1_LVT execution_unit_0_register_file_0_clk_gate_r6_reg (.GCK(
      execution_unit_0_register_file_0_n_65), .CK(cpu_mclk), .E(
      execution_unit_0_register_file_0_n_82), .SE(1'b0));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r6_reg[1] (.Q(
      execution_unit_0_register_file_0_r6[1]), .QN(), .CK(
      execution_unit_0_register_file_0_n_65), .D(
      execution_unit_0_register_file_0_n_67), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_33 (.ZN(
      execution_unit_0_register_file_0_n_105_32), .A1(
      execution_unit_0_register_file_0_n_64), .A2(
      execution_unit_0_register_file_0_r6[1]));
  INV_X1_LVT execution_unit_0_register_file_0_i_27_0 (.ZN(
      execution_unit_0_register_file_0_n_27_0), .A(inst_src[5]));
  NOR2_X1_LVT execution_unit_0_register_file_0_i_27_1 (.ZN(
      execution_unit_0_register_file_0_n_45), .A1(
      execution_unit_0_register_file_0_n_27_0), .A2(execution_unit_0_reg_sr_clr));
  AND2_X1_LVT execution_unit_0_register_file_0_i_29_0 (.ZN(
      execution_unit_0_register_file_0_r5_wr), .A1(inst_dest[5]), .A2(
      execution_unit_0_reg_dest_wr));
  INV_X1_LVT execution_unit_0_register_file_0_i_31_0 (.ZN(
      execution_unit_0_register_file_0_n_31_0), .A(
      execution_unit_0_register_file_0_r5_wr));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_31_3 (.ZN(
      execution_unit_0_register_file_0_n_31_2), .A1(
      execution_unit_0_register_file_0_n_31_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[1]), .B1(
      execution_unit_0_register_file_0_r5_wr), .B2(execution_unit_0_alu_out[1]));
  INV_X1_LVT execution_unit_0_register_file_0_i_31_4 (.ZN(
      execution_unit_0_register_file_0_n_48), .A(
      execution_unit_0_register_file_0_n_31_2));
  AND2_X1_LVT execution_unit_0_register_file_0_i_28_0 (.ZN(
      execution_unit_0_register_file_0_r5_inc), .A1(
      execution_unit_0_register_file_0_n_45), .A2(execution_unit_0_reg_incr));
  INV_X1_LVT execution_unit_0_register_file_0_i_32_1 (.ZN(
      execution_unit_0_register_file_0_n_32_1), .A(
      execution_unit_0_register_file_0_r5_inc));
  INV_X1_LVT execution_unit_0_register_file_0_i_32_0 (.ZN(
      execution_unit_0_register_file_0_n_32_0), .A(
      execution_unit_0_register_file_0_r5_wr));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_32_2 (.ZN(
      execution_unit_0_register_file_0_n_63), .A1(
      execution_unit_0_register_file_0_n_32_1), .A2(
      execution_unit_0_register_file_0_n_32_0));
  CLKGATETST_X1_LVT execution_unit_0_register_file_0_clk_gate_r5_reg (.GCK(
      execution_unit_0_register_file_0_n_46), .CK(cpu_mclk), .E(
      execution_unit_0_register_file_0_n_63), .SE(1'b0));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r5_reg[1] (.Q(
      execution_unit_0_register_file_0_r5[1]), .QN(), .CK(
      execution_unit_0_register_file_0_n_46), .D(
      execution_unit_0_register_file_0_n_48), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_34 (.ZN(
      execution_unit_0_register_file_0_n_105_33), .A1(
      execution_unit_0_register_file_0_n_45), .A2(
      execution_unit_0_register_file_0_r5[1]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_105_35 (.ZN(
      execution_unit_0_register_file_0_n_105_34), .A1(
      execution_unit_0_register_file_0_n_105_30), .A2(
      execution_unit_0_register_file_0_n_105_31), .A3(
      execution_unit_0_register_file_0_n_105_32), .A4(
      execution_unit_0_register_file_0_n_105_33));
  INV_X1_LVT execution_unit_0_register_file_0_i_83_0 (.ZN(
      execution_unit_0_register_file_0_n_83_0), .A(inst_src[13]));
  NOR2_X1_LVT execution_unit_0_register_file_0_i_83_1 (.ZN(
      execution_unit_0_register_file_0_n_197), .A1(
      execution_unit_0_register_file_0_n_83_0), .A2(execution_unit_0_reg_sr_clr));
  AND2_X1_LVT execution_unit_0_register_file_0_i_85_0 (.ZN(
      execution_unit_0_register_file_0_r13_wr), .A1(inst_dest[13]), .A2(
      execution_unit_0_reg_dest_wr));
  INV_X1_LVT execution_unit_0_register_file_0_i_87_0 (.ZN(
      execution_unit_0_register_file_0_n_87_0), .A(
      execution_unit_0_register_file_0_r13_wr));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_87_3 (.ZN(
      execution_unit_0_register_file_0_n_87_2), .A1(
      execution_unit_0_register_file_0_n_87_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[1]), .B1(
      execution_unit_0_register_file_0_r13_wr), .B2(execution_unit_0_alu_out[1]));
  INV_X1_LVT execution_unit_0_register_file_0_i_87_4 (.ZN(
      execution_unit_0_register_file_0_n_200), .A(
      execution_unit_0_register_file_0_n_87_2));
  AND2_X1_LVT execution_unit_0_register_file_0_i_84_0 (.ZN(
      execution_unit_0_register_file_0_r13_inc), .A1(
      execution_unit_0_register_file_0_n_197), .A2(execution_unit_0_reg_incr));
  INV_X1_LVT execution_unit_0_register_file_0_i_88_1 (.ZN(
      execution_unit_0_register_file_0_n_88_1), .A(
      execution_unit_0_register_file_0_r13_inc));
  INV_X1_LVT execution_unit_0_register_file_0_i_88_0 (.ZN(
      execution_unit_0_register_file_0_n_88_0), .A(
      execution_unit_0_register_file_0_r13_wr));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_88_2 (.ZN(
      execution_unit_0_register_file_0_n_215), .A1(
      execution_unit_0_register_file_0_n_88_1), .A2(
      execution_unit_0_register_file_0_n_88_0));
  CLKGATETST_X1_LVT execution_unit_0_register_file_0_clk_gate_r13_reg (.GCK(
      execution_unit_0_register_file_0_n_198), .CK(cpu_mclk), .E(
      execution_unit_0_register_file_0_n_215), .SE(1'b0));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r13_reg[1] (.Q(
      execution_unit_0_register_file_0_r13[1]), .QN(), .CK(
      execution_unit_0_register_file_0_n_198), .D(
      execution_unit_0_register_file_0_n_200), .RN(
      execution_unit_0_register_file_0_n_8));
  AND2_X1_LVT execution_unit_0_register_file_0_i_105_36 (.ZN(
      execution_unit_0_register_file_0_n_105_35), .A1(
      execution_unit_0_register_file_0_n_197), .A2(
      execution_unit_0_register_file_0_r13[1]));
  NOR4_X1_LVT execution_unit_0_register_file_0_i_105_37 (.ZN(
      execution_unit_0_register_file_0_n_105_36), .A1(
      execution_unit_0_register_file_0_n_105_24), .A2(
      execution_unit_0_register_file_0_n_105_29), .A3(
      execution_unit_0_register_file_0_n_105_34), .A4(
      execution_unit_0_register_file_0_n_105_35));
  INV_X1_LVT execution_unit_0_register_file_0_i_104_0 (.ZN(
      execution_unit_0_register_file_0_n_104_0), .A(inst_src[0]));
  NOR2_X1_LVT execution_unit_0_register_file_0_i_104_1 (.ZN(
      execution_unit_0_register_file_0_n_254), .A1(
      execution_unit_0_register_file_0_n_104_0), .A2(execution_unit_0_reg_sr_clr));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_38 (.ZN(
      execution_unit_0_register_file_0_n_105_37), .A1(
      execution_unit_0_register_file_0_n_254), .A2(pc[1]));
  INV_X1_LVT execution_unit_0_register_file_0_i_97_0 (.ZN(
      execution_unit_0_register_file_0_n_97_0), .A(inst_src[15]));
  NOR2_X1_LVT execution_unit_0_register_file_0_i_97_1 (.ZN(
      execution_unit_0_register_file_0_n_235), .A1(
      execution_unit_0_register_file_0_n_97_0), .A2(execution_unit_0_reg_sr_clr));
  AND2_X1_LVT execution_unit_0_register_file_0_i_99_0 (.ZN(
      execution_unit_0_register_file_0_r15_wr), .A1(inst_dest[15]), .A2(
      execution_unit_0_reg_dest_wr));
  INV_X1_LVT execution_unit_0_register_file_0_i_101_0 (.ZN(
      execution_unit_0_register_file_0_n_101_0), .A(
      execution_unit_0_register_file_0_r15_wr));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_101_3 (.ZN(
      execution_unit_0_register_file_0_n_101_2), .A1(
      execution_unit_0_register_file_0_n_101_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[1]), .B1(
      execution_unit_0_register_file_0_r15_wr), .B2(execution_unit_0_alu_out[1]));
  INV_X1_LVT execution_unit_0_register_file_0_i_101_4 (.ZN(
      execution_unit_0_register_file_0_n_238), .A(
      execution_unit_0_register_file_0_n_101_2));
  AND2_X1_LVT execution_unit_0_register_file_0_i_98_0 (.ZN(
      execution_unit_0_register_file_0_r15_inc), .A1(
      execution_unit_0_register_file_0_n_235), .A2(execution_unit_0_reg_incr));
  INV_X1_LVT execution_unit_0_register_file_0_i_102_1 (.ZN(
      execution_unit_0_register_file_0_n_102_1), .A(
      execution_unit_0_register_file_0_r15_inc));
  INV_X1_LVT execution_unit_0_register_file_0_i_102_0 (.ZN(
      execution_unit_0_register_file_0_n_102_0), .A(
      execution_unit_0_register_file_0_r15_wr));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_102_2 (.ZN(
      execution_unit_0_register_file_0_n_253), .A1(
      execution_unit_0_register_file_0_n_102_1), .A2(
      execution_unit_0_register_file_0_n_102_0));
  CLKGATETST_X1_LVT execution_unit_0_register_file_0_clk_gate_r15_reg (.GCK(
      execution_unit_0_register_file_0_n_236), .CK(cpu_mclk), .E(
      execution_unit_0_register_file_0_n_253), .SE(1'b0));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r15_reg[1] (.Q(
      execution_unit_0_register_file_0_r15[1]), .QN(), .CK(
      execution_unit_0_register_file_0_n_236), .D(
      execution_unit_0_register_file_0_n_238), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_39 (.ZN(
      execution_unit_0_register_file_0_n_105_38), .A1(
      execution_unit_0_register_file_0_n_235), .A2(
      execution_unit_0_register_file_0_r15[1]));
  INV_X1_LVT execution_unit_0_register_file_0_i_90_0 (.ZN(
      execution_unit_0_register_file_0_n_90_0), .A(inst_src[14]));
  NOR2_X1_LVT execution_unit_0_register_file_0_i_90_1 (.ZN(
      execution_unit_0_register_file_0_n_216), .A1(
      execution_unit_0_register_file_0_n_90_0), .A2(execution_unit_0_reg_sr_clr));
  AND2_X1_LVT execution_unit_0_register_file_0_i_92_0 (.ZN(
      execution_unit_0_register_file_0_r14_wr), .A1(inst_dest[14]), .A2(
      execution_unit_0_reg_dest_wr));
  INV_X1_LVT execution_unit_0_register_file_0_i_94_0 (.ZN(
      execution_unit_0_register_file_0_n_94_0), .A(
      execution_unit_0_register_file_0_r14_wr));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_94_3 (.ZN(
      execution_unit_0_register_file_0_n_94_2), .A1(
      execution_unit_0_register_file_0_n_94_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[1]), .B1(
      execution_unit_0_register_file_0_r14_wr), .B2(execution_unit_0_alu_out[1]));
  INV_X1_LVT execution_unit_0_register_file_0_i_94_4 (.ZN(
      execution_unit_0_register_file_0_n_219), .A(
      execution_unit_0_register_file_0_n_94_2));
  AND2_X1_LVT execution_unit_0_register_file_0_i_91_0 (.ZN(
      execution_unit_0_register_file_0_r14_inc), .A1(
      execution_unit_0_register_file_0_n_216), .A2(execution_unit_0_reg_incr));
  INV_X1_LVT execution_unit_0_register_file_0_i_95_1 (.ZN(
      execution_unit_0_register_file_0_n_95_1), .A(
      execution_unit_0_register_file_0_r14_inc));
  INV_X1_LVT execution_unit_0_register_file_0_i_95_0 (.ZN(
      execution_unit_0_register_file_0_n_95_0), .A(
      execution_unit_0_register_file_0_r14_wr));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_95_2 (.ZN(
      execution_unit_0_register_file_0_n_234), .A1(
      execution_unit_0_register_file_0_n_95_1), .A2(
      execution_unit_0_register_file_0_n_95_0));
  CLKGATETST_X1_LVT execution_unit_0_register_file_0_clk_gate_r14_reg (.GCK(
      execution_unit_0_register_file_0_n_217), .CK(cpu_mclk), .E(
      execution_unit_0_register_file_0_n_234), .SE(1'b0));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r14_reg[1] (.Q(
      execution_unit_0_register_file_0_r14[1]), .QN(), .CK(
      execution_unit_0_register_file_0_n_217), .D(
      execution_unit_0_register_file_0_n_219), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_40 (.ZN(
      execution_unit_0_register_file_0_n_105_39), .A1(
      execution_unit_0_register_file_0_n_216), .A2(
      execution_unit_0_register_file_0_r14[1]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_105_41 (.ZN(
      execution_unit_0_reg_src[1]), .A1(
      execution_unit_0_register_file_0_n_105_36), .A2(
      execution_unit_0_register_file_0_n_105_37), .A3(
      execution_unit_0_register_file_0_n_105_38), .A4(
      execution_unit_0_register_file_0_n_105_39));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_24_1 (.ZN(
      execution_unit_0_register_file_0_n_24_1), .A1(
      execution_unit_0_register_file_0_n_24_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[0]), .B1(
      execution_unit_0_alu_out[0]), .B2(execution_unit_0_register_file_0_r4_wr));
  INV_X1_LVT execution_unit_0_register_file_0_i_24_2 (.ZN(
      execution_unit_0_register_file_0_n_28), .A(
      execution_unit_0_register_file_0_n_24_1));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r4_reg[0] (.Q(
      execution_unit_0_register_file_0_r4[0]), .QN(), .CK(
      execution_unit_0_register_file_0_n_27), .D(
      execution_unit_0_register_file_0_n_28), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_0 (.ZN(
      execution_unit_0_register_file_0_n_105_0), .A1(
      execution_unit_0_register_file_0_r4[0]), .A2(
      execution_unit_0_register_file_0_n_24));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r3_reg[0] (.Q(
      execution_unit_0_register_file_0_r3[0]), .QN(), .CK(
      execution_unit_0_register_file_0_n_23), .D(execution_unit_0_alu_out[0]), 
      .RN(execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_1 (.ZN(
      execution_unit_0_register_file_0_n_105_1), .A1(
      execution_unit_0_register_file_0_r3[0]), .A2(
      execution_unit_0_register_file_0_n_22));
  INV_X1_LVT execution_unit_0_register_file_0_i_5_1 (.ZN(
      execution_unit_0_register_file_0_n_5_1), .A(execution_unit_0_alu_stat_wr[0]));
  NAND3_X1_LVT execution_unit_0_register_file_0_i_5_2 (.ZN(
      execution_unit_0_register_file_0_n_5_2), .A1(
      execution_unit_0_register_file_0_n_5_0), .A2(
      execution_unit_0_register_file_0_n_5_1), .A3(execution_unit_0_status[0]));
  NAND3_X1_LVT execution_unit_0_register_file_0_i_5_3 (.ZN(
      execution_unit_0_register_file_0_n_5_3), .A1(
      execution_unit_0_register_file_0_n_5_1), .A2(
      execution_unit_0_register_file_0_r2_wr), .A3(execution_unit_0_alu_out[0]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_5_4 (.ZN(
      execution_unit_0_register_file_0_n_5_4), .A1(execution_unit_0_alu_stat[0]), 
      .A2(execution_unit_0_alu_stat_wr[0]));
  NAND3_X1_LVT execution_unit_0_register_file_0_i_5_5 (.ZN(
      execution_unit_0_register_file_0_n_9), .A1(
      execution_unit_0_register_file_0_n_5_2), .A2(
      execution_unit_0_register_file_0_n_5_3), .A3(
      execution_unit_0_register_file_0_n_5_4));
  AND2_X1_LVT execution_unit_0_register_file_0_i_6_1 (.ZN(
      execution_unit_0_register_file_0_n_13), .A1(
      execution_unit_0_register_file_0_n_6_0), .A2(
      execution_unit_0_register_file_0_n_9));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r2_reg[0] (.Q(
      execution_unit_0_status[0]), .QN(), .CK(cpu_mclk), .D(
      execution_unit_0_register_file_0_n_13), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_2 (.ZN(
      execution_unit_0_register_file_0_n_105_2), .A1(execution_unit_0_status[0]), 
      .A2(execution_unit_0_register_file_0_n_21));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r1_reg[0] (.Q(
      execution_unit_0_register_file_0_r1[0]), .QN(), .CK(
      execution_unit_0_register_file_0_n_270), .D(1'b0), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_3 (.ZN(
      execution_unit_0_register_file_0_n_105_3), .A1(
      execution_unit_0_register_file_0_r1[0]), .A2(
      execution_unit_0_register_file_0_inst_src_in));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_105_4 (.ZN(
      execution_unit_0_register_file_0_n_105_4), .A1(
      execution_unit_0_register_file_0_n_105_0), .A2(
      execution_unit_0_register_file_0_n_105_1), .A3(
      execution_unit_0_register_file_0_n_105_2), .A4(
      execution_unit_0_register_file_0_n_105_3));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_80_1 (.ZN(
      execution_unit_0_register_file_0_n_80_1), .A1(
      execution_unit_0_register_file_0_n_80_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[0]), .B1(
      execution_unit_0_alu_out[0]), .B2(execution_unit_0_register_file_0_r12_wr));
  INV_X1_LVT execution_unit_0_register_file_0_i_80_2 (.ZN(
      execution_unit_0_register_file_0_n_180), .A(
      execution_unit_0_register_file_0_n_80_1));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r12_reg[0] (.Q(
      execution_unit_0_register_file_0_r12[0]), .QN(), .CK(
      execution_unit_0_register_file_0_n_179), .D(
      execution_unit_0_register_file_0_n_180), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_5 (.ZN(
      execution_unit_0_register_file_0_n_105_5), .A1(
      execution_unit_0_register_file_0_r12[0]), .A2(
      execution_unit_0_register_file_0_n_178));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_73_1 (.ZN(
      execution_unit_0_register_file_0_n_73_1), .A1(
      execution_unit_0_register_file_0_n_73_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[0]), .B1(
      execution_unit_0_alu_out[0]), .B2(execution_unit_0_register_file_0_r11_wr));
  INV_X1_LVT execution_unit_0_register_file_0_i_73_2 (.ZN(
      execution_unit_0_register_file_0_n_161), .A(
      execution_unit_0_register_file_0_n_73_1));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r11_reg[0] (.Q(
      execution_unit_0_register_file_0_r11[0]), .QN(), .CK(
      execution_unit_0_register_file_0_n_160), .D(
      execution_unit_0_register_file_0_n_161), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_6 (.ZN(
      execution_unit_0_register_file_0_n_105_6), .A1(
      execution_unit_0_register_file_0_r11[0]), .A2(
      execution_unit_0_register_file_0_n_159));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_66_1 (.ZN(
      execution_unit_0_register_file_0_n_66_1), .A1(
      execution_unit_0_register_file_0_n_66_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[0]), .B1(
      execution_unit_0_alu_out[0]), .B2(execution_unit_0_register_file_0_r10_wr));
  INV_X1_LVT execution_unit_0_register_file_0_i_66_2 (.ZN(
      execution_unit_0_register_file_0_n_142), .A(
      execution_unit_0_register_file_0_n_66_1));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r10_reg[0] (.Q(
      execution_unit_0_register_file_0_r10[0]), .QN(), .CK(
      execution_unit_0_register_file_0_n_141), .D(
      execution_unit_0_register_file_0_n_142), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_7 (.ZN(
      execution_unit_0_register_file_0_n_105_7), .A1(
      execution_unit_0_register_file_0_r10[0]), .A2(
      execution_unit_0_register_file_0_n_140));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_59_1 (.ZN(
      execution_unit_0_register_file_0_n_59_1), .A1(
      execution_unit_0_register_file_0_n_59_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[0]), .B1(
      execution_unit_0_alu_out[0]), .B2(execution_unit_0_register_file_0_r9_wr));
  INV_X1_LVT execution_unit_0_register_file_0_i_59_2 (.ZN(
      execution_unit_0_register_file_0_n_123), .A(
      execution_unit_0_register_file_0_n_59_1));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r9_reg[0] (.Q(
      execution_unit_0_register_file_0_r9[0]), .QN(), .CK(
      execution_unit_0_register_file_0_n_122), .D(
      execution_unit_0_register_file_0_n_123), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_8 (.ZN(
      execution_unit_0_register_file_0_n_105_8), .A1(
      execution_unit_0_register_file_0_r9[0]), .A2(
      execution_unit_0_register_file_0_n_121));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_105_9 (.ZN(
      execution_unit_0_register_file_0_n_105_9), .A1(
      execution_unit_0_register_file_0_n_105_5), .A2(
      execution_unit_0_register_file_0_n_105_6), .A3(
      execution_unit_0_register_file_0_n_105_7), .A4(
      execution_unit_0_register_file_0_n_105_8));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_52_1 (.ZN(
      execution_unit_0_register_file_0_n_52_1), .A1(
      execution_unit_0_register_file_0_n_52_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[0]), .B1(
      execution_unit_0_alu_out[0]), .B2(execution_unit_0_register_file_0_r8_wr));
  INV_X1_LVT execution_unit_0_register_file_0_i_52_2 (.ZN(
      execution_unit_0_register_file_0_n_104), .A(
      execution_unit_0_register_file_0_n_52_1));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r8_reg[0] (.Q(
      execution_unit_0_register_file_0_r8[0]), .QN(), .CK(
      execution_unit_0_register_file_0_n_103), .D(
      execution_unit_0_register_file_0_n_104), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_10 (.ZN(
      execution_unit_0_register_file_0_n_105_10), .A1(
      execution_unit_0_register_file_0_r8[0]), .A2(
      execution_unit_0_register_file_0_n_102));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_45_1 (.ZN(
      execution_unit_0_register_file_0_n_45_1), .A1(
      execution_unit_0_register_file_0_n_45_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[0]), .B1(
      execution_unit_0_alu_out[0]), .B2(execution_unit_0_register_file_0_r7_wr));
  INV_X1_LVT execution_unit_0_register_file_0_i_45_2 (.ZN(
      execution_unit_0_register_file_0_n_85), .A(
      execution_unit_0_register_file_0_n_45_1));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r7_reg[0] (.Q(
      execution_unit_0_register_file_0_r7[0]), .QN(), .CK(
      execution_unit_0_register_file_0_n_84), .D(
      execution_unit_0_register_file_0_n_85), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_11 (.ZN(
      execution_unit_0_register_file_0_n_105_11), .A1(
      execution_unit_0_register_file_0_r7[0]), .A2(
      execution_unit_0_register_file_0_n_83));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_38_1 (.ZN(
      execution_unit_0_register_file_0_n_38_1), .A1(
      execution_unit_0_register_file_0_n_38_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[0]), .B1(
      execution_unit_0_alu_out[0]), .B2(execution_unit_0_register_file_0_r6_wr));
  INV_X1_LVT execution_unit_0_register_file_0_i_38_2 (.ZN(
      execution_unit_0_register_file_0_n_66), .A(
      execution_unit_0_register_file_0_n_38_1));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r6_reg[0] (.Q(
      execution_unit_0_register_file_0_r6[0]), .QN(), .CK(
      execution_unit_0_register_file_0_n_65), .D(
      execution_unit_0_register_file_0_n_66), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_12 (.ZN(
      execution_unit_0_register_file_0_n_105_12), .A1(
      execution_unit_0_register_file_0_r6[0]), .A2(
      execution_unit_0_register_file_0_n_64));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_31_1 (.ZN(
      execution_unit_0_register_file_0_n_31_1), .A1(
      execution_unit_0_register_file_0_n_31_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[0]), .B1(
      execution_unit_0_alu_out[0]), .B2(execution_unit_0_register_file_0_r5_wr));
  INV_X1_LVT execution_unit_0_register_file_0_i_31_2 (.ZN(
      execution_unit_0_register_file_0_n_47), .A(
      execution_unit_0_register_file_0_n_31_1));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r5_reg[0] (.Q(
      execution_unit_0_register_file_0_r5[0]), .QN(), .CK(
      execution_unit_0_register_file_0_n_46), .D(
      execution_unit_0_register_file_0_n_47), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_13 (.ZN(
      execution_unit_0_register_file_0_n_105_13), .A1(
      execution_unit_0_register_file_0_r5[0]), .A2(
      execution_unit_0_register_file_0_n_45));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_105_14 (.ZN(
      execution_unit_0_register_file_0_n_105_14), .A1(
      execution_unit_0_register_file_0_n_105_10), .A2(
      execution_unit_0_register_file_0_n_105_11), .A3(
      execution_unit_0_register_file_0_n_105_12), .A4(
      execution_unit_0_register_file_0_n_105_13));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_87_1 (.ZN(
      execution_unit_0_register_file_0_n_87_1), .A1(
      execution_unit_0_register_file_0_n_87_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[0]), .B1(
      execution_unit_0_alu_out[0]), .B2(execution_unit_0_register_file_0_r13_wr));
  INV_X1_LVT execution_unit_0_register_file_0_i_87_2 (.ZN(
      execution_unit_0_register_file_0_n_199), .A(
      execution_unit_0_register_file_0_n_87_1));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r13_reg[0] (.Q(
      execution_unit_0_register_file_0_r13[0]), .QN(), .CK(
      execution_unit_0_register_file_0_n_198), .D(
      execution_unit_0_register_file_0_n_199), .RN(
      execution_unit_0_register_file_0_n_8));
  AND2_X1_LVT execution_unit_0_register_file_0_i_105_15 (.ZN(
      execution_unit_0_register_file_0_n_105_15), .A1(
      execution_unit_0_register_file_0_r13[0]), .A2(
      execution_unit_0_register_file_0_n_197));
  NOR4_X1_LVT execution_unit_0_register_file_0_i_105_16 (.ZN(
      execution_unit_0_register_file_0_n_105_16), .A1(
      execution_unit_0_register_file_0_n_105_4), .A2(
      execution_unit_0_register_file_0_n_105_9), .A3(
      execution_unit_0_register_file_0_n_105_14), .A4(
      execution_unit_0_register_file_0_n_105_15));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_17 (.ZN(
      execution_unit_0_register_file_0_n_105_17), .A1(pc[0]), .A2(
      execution_unit_0_register_file_0_n_254));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_101_1 (.ZN(
      execution_unit_0_register_file_0_n_101_1), .A1(
      execution_unit_0_register_file_0_n_101_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[0]), .B1(
      execution_unit_0_alu_out[0]), .B2(execution_unit_0_register_file_0_r15_wr));
  INV_X1_LVT execution_unit_0_register_file_0_i_101_2 (.ZN(
      execution_unit_0_register_file_0_n_237), .A(
      execution_unit_0_register_file_0_n_101_1));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r15_reg[0] (.Q(
      execution_unit_0_register_file_0_r15[0]), .QN(), .CK(
      execution_unit_0_register_file_0_n_236), .D(
      execution_unit_0_register_file_0_n_237), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_18 (.ZN(
      execution_unit_0_register_file_0_n_105_18), .A1(
      execution_unit_0_register_file_0_r15[0]), .A2(
      execution_unit_0_register_file_0_n_235));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_94_1 (.ZN(
      execution_unit_0_register_file_0_n_94_1), .A1(
      execution_unit_0_register_file_0_n_94_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[0]), .B1(
      execution_unit_0_alu_out[0]), .B2(execution_unit_0_register_file_0_r14_wr));
  INV_X1_LVT execution_unit_0_register_file_0_i_94_2 (.ZN(
      execution_unit_0_register_file_0_n_218), .A(
      execution_unit_0_register_file_0_n_94_1));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r14_reg[0] (.Q(
      execution_unit_0_register_file_0_r14[0]), .QN(), .CK(
      execution_unit_0_register_file_0_n_217), .D(
      execution_unit_0_register_file_0_n_218), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_19 (.ZN(
      execution_unit_0_register_file_0_n_105_19), .A1(
      execution_unit_0_register_file_0_r14[0]), .A2(
      execution_unit_0_register_file_0_n_216));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_105_20 (.ZN(
      execution_unit_0_reg_src[0]), .A1(execution_unit_0_register_file_0_n_105_16), 
      .A2(execution_unit_0_register_file_0_n_105_17), .A3(
      execution_unit_0_register_file_0_n_105_18), .A4(
      execution_unit_0_register_file_0_n_105_19));
  HA_X1_LVT execution_unit_0_register_file_0_i_22_0 (.CO(
      execution_unit_0_register_file_0_n_22_0), .S(
      execution_unit_0_register_file_0_reg_incr_val[0]), .A(
      execution_unit_0_register_file_0_n_25), .B(execution_unit_0_reg_src[0]));
  FA_X1_LVT execution_unit_0_register_file_0_i_22_1 (.CO(
      execution_unit_0_register_file_0_n_22_1), .S(
      execution_unit_0_register_file_0_reg_incr_val[1]), .A(
      execution_unit_0_register_file_0_n_26), .B(execution_unit_0_reg_src[1]), 
      .CI(execution_unit_0_register_file_0_n_22_0));
  HA_X1_LVT execution_unit_0_register_file_0_i_22_2 (.CO(
      execution_unit_0_register_file_0_n_22_2), .S(
      execution_unit_0_register_file_0_reg_incr_val[2]), .A(
      execution_unit_0_reg_src[2]), .B(execution_unit_0_register_file_0_n_22_1));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_24_5 (.ZN(
      execution_unit_0_register_file_0_n_24_3), .A1(
      execution_unit_0_register_file_0_n_24_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[2]), .B1(
      execution_unit_0_register_file_0_r4_wr), .B2(execution_unit_0_alu_out[2]));
  INV_X1_LVT execution_unit_0_register_file_0_i_24_6 (.ZN(
      execution_unit_0_register_file_0_n_30), .A(
      execution_unit_0_register_file_0_n_24_3));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r4_reg[2] (.Q(
      execution_unit_0_register_file_0_r4[2]), .QN(), .CK(
      execution_unit_0_register_file_0_n_27), .D(
      execution_unit_0_register_file_0_n_30), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_42 (.ZN(
      execution_unit_0_register_file_0_n_105_40), .A1(
      execution_unit_0_register_file_0_n_24), .A2(
      execution_unit_0_register_file_0_r4[2]));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r3_reg[2] (.Q(
      execution_unit_0_register_file_0_r3[2]), .QN(), .CK(
      execution_unit_0_register_file_0_n_23), .D(execution_unit_0_alu_out[2]), 
      .RN(execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_43 (.ZN(
      execution_unit_0_register_file_0_n_105_41), .A1(
      execution_unit_0_register_file_0_n_22), .A2(
      execution_unit_0_register_file_0_r3[2]));
  INV_X1_LVT execution_unit_0_register_file_0_i_5_11 (.ZN(
      execution_unit_0_register_file_0_n_5_9), .A(
      execution_unit_0_alu_stat_wr[2]));
  NAND3_X1_LVT execution_unit_0_register_file_0_i_5_12 (.ZN(
      execution_unit_0_register_file_0_n_5_10), .A1(
      execution_unit_0_register_file_0_n_5_0), .A2(
      execution_unit_0_register_file_0_n_5_9), .A3(execution_unit_0_status[2]));
  NAND3_X1_LVT execution_unit_0_register_file_0_i_5_13 (.ZN(
      execution_unit_0_register_file_0_n_5_11), .A1(
      execution_unit_0_register_file_0_n_5_9), .A2(
      execution_unit_0_register_file_0_r2_wr), .A3(execution_unit_0_alu_out[2]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_5_14 (.ZN(
      execution_unit_0_register_file_0_n_5_12), .A1(execution_unit_0_alu_stat[2]), 
      .A2(execution_unit_0_alu_stat_wr[2]));
  NAND3_X1_LVT execution_unit_0_register_file_0_i_5_15 (.ZN(
      execution_unit_0_register_file_0_n_11), .A1(
      execution_unit_0_register_file_0_n_5_10), .A2(
      execution_unit_0_register_file_0_n_5_11), .A3(
      execution_unit_0_register_file_0_n_5_12));
  AND2_X1_LVT execution_unit_0_register_file_0_i_6_3 (.ZN(
      execution_unit_0_register_file_0_n_15), .A1(
      execution_unit_0_register_file_0_n_6_0), .A2(
      execution_unit_0_register_file_0_n_11));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r2_reg[2] (.Q(
      execution_unit_0_status[2]), .QN(), .CK(cpu_mclk), .D(
      execution_unit_0_register_file_0_n_15), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_44 (.ZN(
      execution_unit_0_register_file_0_n_105_42), .A1(
      execution_unit_0_register_file_0_n_21), .A2(execution_unit_0_status[2]));
  AOI222_X1_LVT execution_unit_0_register_file_0_i_109_2 (.ZN(
      execution_unit_0_register_file_0_n_109_1), .A1(
      execution_unit_0_register_file_0_r1_wr), .A2(execution_unit_0_alu_out[2]), 
      .B1(execution_unit_0_register_file_0_n_272), .B2(eu_mab[2]), .C1(
      execution_unit_0_register_file_0_n_271), .C2(
      execution_unit_0_register_file_0_n_256));
  INV_X1_LVT execution_unit_0_register_file_0_i_109_3 (.ZN(
      execution_unit_0_register_file_0_n_274), .A(
      execution_unit_0_register_file_0_n_109_1));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r1_reg[2] (.Q(
      execution_unit_0_register_file_0_r1[2]), .QN(), .CK(
      execution_unit_0_register_file_0_n_270), .D(
      execution_unit_0_register_file_0_n_274), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_45 (.ZN(
      execution_unit_0_register_file_0_n_105_43), .A1(
      execution_unit_0_register_file_0_inst_src_in), .A2(
      execution_unit_0_register_file_0_r1[2]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_105_46 (.ZN(
      execution_unit_0_register_file_0_n_105_44), .A1(
      execution_unit_0_register_file_0_n_105_40), .A2(
      execution_unit_0_register_file_0_n_105_41), .A3(
      execution_unit_0_register_file_0_n_105_42), .A4(
      execution_unit_0_register_file_0_n_105_43));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_80_5 (.ZN(
      execution_unit_0_register_file_0_n_80_3), .A1(
      execution_unit_0_register_file_0_n_80_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[2]), .B1(
      execution_unit_0_register_file_0_r12_wr), .B2(execution_unit_0_alu_out[2]));
  INV_X1_LVT execution_unit_0_register_file_0_i_80_6 (.ZN(
      execution_unit_0_register_file_0_n_182), .A(
      execution_unit_0_register_file_0_n_80_3));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r12_reg[2] (.Q(
      execution_unit_0_register_file_0_r12[2]), .QN(), .CK(
      execution_unit_0_register_file_0_n_179), .D(
      execution_unit_0_register_file_0_n_182), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_47 (.ZN(
      execution_unit_0_register_file_0_n_105_45), .A1(
      execution_unit_0_register_file_0_n_178), .A2(
      execution_unit_0_register_file_0_r12[2]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_73_5 (.ZN(
      execution_unit_0_register_file_0_n_73_3), .A1(
      execution_unit_0_register_file_0_n_73_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[2]), .B1(
      execution_unit_0_register_file_0_r11_wr), .B2(execution_unit_0_alu_out[2]));
  INV_X1_LVT execution_unit_0_register_file_0_i_73_6 (.ZN(
      execution_unit_0_register_file_0_n_163), .A(
      execution_unit_0_register_file_0_n_73_3));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r11_reg[2] (.Q(
      execution_unit_0_register_file_0_r11[2]), .QN(), .CK(
      execution_unit_0_register_file_0_n_160), .D(
      execution_unit_0_register_file_0_n_163), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_48 (.ZN(
      execution_unit_0_register_file_0_n_105_46), .A1(
      execution_unit_0_register_file_0_n_159), .A2(
      execution_unit_0_register_file_0_r11[2]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_66_5 (.ZN(
      execution_unit_0_register_file_0_n_66_3), .A1(
      execution_unit_0_register_file_0_n_66_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[2]), .B1(
      execution_unit_0_register_file_0_r10_wr), .B2(execution_unit_0_alu_out[2]));
  INV_X1_LVT execution_unit_0_register_file_0_i_66_6 (.ZN(
      execution_unit_0_register_file_0_n_144), .A(
      execution_unit_0_register_file_0_n_66_3));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r10_reg[2] (.Q(
      execution_unit_0_register_file_0_r10[2]), .QN(), .CK(
      execution_unit_0_register_file_0_n_141), .D(
      execution_unit_0_register_file_0_n_144), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_49 (.ZN(
      execution_unit_0_register_file_0_n_105_47), .A1(
      execution_unit_0_register_file_0_n_140), .A2(
      execution_unit_0_register_file_0_r10[2]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_59_5 (.ZN(
      execution_unit_0_register_file_0_n_59_3), .A1(
      execution_unit_0_register_file_0_n_59_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[2]), .B1(
      execution_unit_0_register_file_0_r9_wr), .B2(execution_unit_0_alu_out[2]));
  INV_X1_LVT execution_unit_0_register_file_0_i_59_6 (.ZN(
      execution_unit_0_register_file_0_n_125), .A(
      execution_unit_0_register_file_0_n_59_3));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r9_reg[2] (.Q(
      execution_unit_0_register_file_0_r9[2]), .QN(), .CK(
      execution_unit_0_register_file_0_n_122), .D(
      execution_unit_0_register_file_0_n_125), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_50 (.ZN(
      execution_unit_0_register_file_0_n_105_48), .A1(
      execution_unit_0_register_file_0_n_121), .A2(
      execution_unit_0_register_file_0_r9[2]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_105_51 (.ZN(
      execution_unit_0_register_file_0_n_105_49), .A1(
      execution_unit_0_register_file_0_n_105_45), .A2(
      execution_unit_0_register_file_0_n_105_46), .A3(
      execution_unit_0_register_file_0_n_105_47), .A4(
      execution_unit_0_register_file_0_n_105_48));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_52_5 (.ZN(
      execution_unit_0_register_file_0_n_52_3), .A1(
      execution_unit_0_register_file_0_n_52_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[2]), .B1(
      execution_unit_0_register_file_0_r8_wr), .B2(execution_unit_0_alu_out[2]));
  INV_X1_LVT execution_unit_0_register_file_0_i_52_6 (.ZN(
      execution_unit_0_register_file_0_n_106), .A(
      execution_unit_0_register_file_0_n_52_3));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r8_reg[2] (.Q(
      execution_unit_0_register_file_0_r8[2]), .QN(), .CK(
      execution_unit_0_register_file_0_n_103), .D(
      execution_unit_0_register_file_0_n_106), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_52 (.ZN(
      execution_unit_0_register_file_0_n_105_50), .A1(
      execution_unit_0_register_file_0_n_102), .A2(
      execution_unit_0_register_file_0_r8[2]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_45_5 (.ZN(
      execution_unit_0_register_file_0_n_45_3), .A1(
      execution_unit_0_register_file_0_n_45_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[2]), .B1(
      execution_unit_0_register_file_0_r7_wr), .B2(execution_unit_0_alu_out[2]));
  INV_X1_LVT execution_unit_0_register_file_0_i_45_6 (.ZN(
      execution_unit_0_register_file_0_n_87), .A(
      execution_unit_0_register_file_0_n_45_3));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r7_reg[2] (.Q(
      execution_unit_0_register_file_0_r7[2]), .QN(), .CK(
      execution_unit_0_register_file_0_n_84), .D(
      execution_unit_0_register_file_0_n_87), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_53 (.ZN(
      execution_unit_0_register_file_0_n_105_51), .A1(
      execution_unit_0_register_file_0_n_83), .A2(
      execution_unit_0_register_file_0_r7[2]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_38_5 (.ZN(
      execution_unit_0_register_file_0_n_38_3), .A1(
      execution_unit_0_register_file_0_n_38_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[2]), .B1(
      execution_unit_0_register_file_0_r6_wr), .B2(execution_unit_0_alu_out[2]));
  INV_X1_LVT execution_unit_0_register_file_0_i_38_6 (.ZN(
      execution_unit_0_register_file_0_n_68), .A(
      execution_unit_0_register_file_0_n_38_3));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r6_reg[2] (.Q(
      execution_unit_0_register_file_0_r6[2]), .QN(), .CK(
      execution_unit_0_register_file_0_n_65), .D(
      execution_unit_0_register_file_0_n_68), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_54 (.ZN(
      execution_unit_0_register_file_0_n_105_52), .A1(
      execution_unit_0_register_file_0_n_64), .A2(
      execution_unit_0_register_file_0_r6[2]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_31_5 (.ZN(
      execution_unit_0_register_file_0_n_31_3), .A1(
      execution_unit_0_register_file_0_n_31_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[2]), .B1(
      execution_unit_0_register_file_0_r5_wr), .B2(execution_unit_0_alu_out[2]));
  INV_X1_LVT execution_unit_0_register_file_0_i_31_6 (.ZN(
      execution_unit_0_register_file_0_n_49), .A(
      execution_unit_0_register_file_0_n_31_3));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r5_reg[2] (.Q(
      execution_unit_0_register_file_0_r5[2]), .QN(), .CK(
      execution_unit_0_register_file_0_n_46), .D(
      execution_unit_0_register_file_0_n_49), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_55 (.ZN(
      execution_unit_0_register_file_0_n_105_53), .A1(
      execution_unit_0_register_file_0_n_45), .A2(
      execution_unit_0_register_file_0_r5[2]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_105_56 (.ZN(
      execution_unit_0_register_file_0_n_105_54), .A1(
      execution_unit_0_register_file_0_n_105_50), .A2(
      execution_unit_0_register_file_0_n_105_51), .A3(
      execution_unit_0_register_file_0_n_105_52), .A4(
      execution_unit_0_register_file_0_n_105_53));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_87_5 (.ZN(
      execution_unit_0_register_file_0_n_87_3), .A1(
      execution_unit_0_register_file_0_n_87_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[2]), .B1(
      execution_unit_0_register_file_0_r13_wr), .B2(execution_unit_0_alu_out[2]));
  INV_X1_LVT execution_unit_0_register_file_0_i_87_6 (.ZN(
      execution_unit_0_register_file_0_n_201), .A(
      execution_unit_0_register_file_0_n_87_3));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r13_reg[2] (.Q(
      execution_unit_0_register_file_0_r13[2]), .QN(), .CK(
      execution_unit_0_register_file_0_n_198), .D(
      execution_unit_0_register_file_0_n_201), .RN(
      execution_unit_0_register_file_0_n_8));
  AND2_X1_LVT execution_unit_0_register_file_0_i_105_57 (.ZN(
      execution_unit_0_register_file_0_n_105_55), .A1(
      execution_unit_0_register_file_0_n_197), .A2(
      execution_unit_0_register_file_0_r13[2]));
  NOR4_X1_LVT execution_unit_0_register_file_0_i_105_58 (.ZN(
      execution_unit_0_register_file_0_n_105_56), .A1(
      execution_unit_0_register_file_0_n_105_44), .A2(
      execution_unit_0_register_file_0_n_105_49), .A3(
      execution_unit_0_register_file_0_n_105_54), .A4(
      execution_unit_0_register_file_0_n_105_55));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_59 (.ZN(
      execution_unit_0_register_file_0_n_105_57), .A1(
      execution_unit_0_register_file_0_n_254), .A2(pc[2]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_101_5 (.ZN(
      execution_unit_0_register_file_0_n_101_3), .A1(
      execution_unit_0_register_file_0_n_101_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[2]), .B1(
      execution_unit_0_register_file_0_r15_wr), .B2(execution_unit_0_alu_out[2]));
  INV_X1_LVT execution_unit_0_register_file_0_i_101_6 (.ZN(
      execution_unit_0_register_file_0_n_239), .A(
      execution_unit_0_register_file_0_n_101_3));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r15_reg[2] (.Q(
      execution_unit_0_register_file_0_r15[2]), .QN(), .CK(
      execution_unit_0_register_file_0_n_236), .D(
      execution_unit_0_register_file_0_n_239), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_60 (.ZN(
      execution_unit_0_register_file_0_n_105_58), .A1(
      execution_unit_0_register_file_0_n_235), .A2(
      execution_unit_0_register_file_0_r15[2]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_94_5 (.ZN(
      execution_unit_0_register_file_0_n_94_3), .A1(
      execution_unit_0_register_file_0_n_94_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[2]), .B1(
      execution_unit_0_register_file_0_r14_wr), .B2(execution_unit_0_alu_out[2]));
  INV_X1_LVT execution_unit_0_register_file_0_i_94_6 (.ZN(
      execution_unit_0_register_file_0_n_220), .A(
      execution_unit_0_register_file_0_n_94_3));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r14_reg[2] (.Q(
      execution_unit_0_register_file_0_r14[2]), .QN(), .CK(
      execution_unit_0_register_file_0_n_217), .D(
      execution_unit_0_register_file_0_n_220), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_61 (.ZN(
      execution_unit_0_register_file_0_n_105_59), .A1(
      execution_unit_0_register_file_0_n_216), .A2(
      execution_unit_0_register_file_0_r14[2]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_105_62 (.ZN(
      execution_unit_0_reg_src[2]), .A1(
      execution_unit_0_register_file_0_n_105_56), .A2(
      execution_unit_0_register_file_0_n_105_57), .A3(
      execution_unit_0_register_file_0_n_105_58), .A4(
      execution_unit_0_register_file_0_n_105_59));
  HA_X1_LVT execution_unit_0_register_file_0_i_106_1 (.CO(
      execution_unit_0_register_file_0_n_106_0), .S(
      execution_unit_0_register_file_0_n_256), .A(execution_unit_0_reg_src[2]), 
      .B(execution_unit_0_reg_src[1]));
  HA_X1_LVT execution_unit_0_register_file_0_i_106_2 (.CO(
      execution_unit_0_register_file_0_n_106_1), .S(
      execution_unit_0_register_file_0_n_257), .A(execution_unit_0_reg_src[3]), 
      .B(execution_unit_0_register_file_0_n_106_0));
  AOI222_X1_LVT execution_unit_0_register_file_0_i_109_4 (.ZN(
      execution_unit_0_register_file_0_n_109_2), .A1(
      execution_unit_0_register_file_0_r1_wr), .A2(execution_unit_0_alu_out[3]), 
      .B1(execution_unit_0_register_file_0_n_272), .B2(eu_mab[3]), .C1(
      execution_unit_0_register_file_0_n_271), .C2(
      execution_unit_0_register_file_0_n_257));
  INV_X1_LVT execution_unit_0_register_file_0_i_109_5 (.ZN(
      execution_unit_0_register_file_0_n_275), .A(
      execution_unit_0_register_file_0_n_109_2));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r1_reg[3] (.Q(
      execution_unit_0_register_file_0_r1[3]), .QN(), .CK(
      execution_unit_0_register_file_0_n_270), .D(
      execution_unit_0_register_file_0_n_275), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_66 (.ZN(
      execution_unit_0_register_file_0_n_105_63), .A1(
      execution_unit_0_register_file_0_inst_src_in), .A2(
      execution_unit_0_register_file_0_r1[3]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_105_67 (.ZN(
      execution_unit_0_register_file_0_n_105_64), .A1(
      execution_unit_0_register_file_0_n_105_60), .A2(
      execution_unit_0_register_file_0_n_105_61), .A3(
      execution_unit_0_register_file_0_n_105_62), .A4(
      execution_unit_0_register_file_0_n_105_63));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_80_7 (.ZN(
      execution_unit_0_register_file_0_n_80_4), .A1(
      execution_unit_0_register_file_0_n_80_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[3]), .B1(
      execution_unit_0_register_file_0_r12_wr), .B2(execution_unit_0_alu_out[3]));
  INV_X1_LVT execution_unit_0_register_file_0_i_80_8 (.ZN(
      execution_unit_0_register_file_0_n_183), .A(
      execution_unit_0_register_file_0_n_80_4));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r12_reg[3] (.Q(
      execution_unit_0_register_file_0_r12[3]), .QN(), .CK(
      execution_unit_0_register_file_0_n_179), .D(
      execution_unit_0_register_file_0_n_183), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_68 (.ZN(
      execution_unit_0_register_file_0_n_105_65), .A1(
      execution_unit_0_register_file_0_n_178), .A2(
      execution_unit_0_register_file_0_r12[3]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_73_7 (.ZN(
      execution_unit_0_register_file_0_n_73_4), .A1(
      execution_unit_0_register_file_0_n_73_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[3]), .B1(
      execution_unit_0_register_file_0_r11_wr), .B2(execution_unit_0_alu_out[3]));
  INV_X1_LVT execution_unit_0_register_file_0_i_73_8 (.ZN(
      execution_unit_0_register_file_0_n_164), .A(
      execution_unit_0_register_file_0_n_73_4));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r11_reg[3] (.Q(
      execution_unit_0_register_file_0_r11[3]), .QN(), .CK(
      execution_unit_0_register_file_0_n_160), .D(
      execution_unit_0_register_file_0_n_164), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_69 (.ZN(
      execution_unit_0_register_file_0_n_105_66), .A1(
      execution_unit_0_register_file_0_n_159), .A2(
      execution_unit_0_register_file_0_r11[3]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_66_7 (.ZN(
      execution_unit_0_register_file_0_n_66_4), .A1(
      execution_unit_0_register_file_0_n_66_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[3]), .B1(
      execution_unit_0_register_file_0_r10_wr), .B2(execution_unit_0_alu_out[3]));
  INV_X1_LVT execution_unit_0_register_file_0_i_66_8 (.ZN(
      execution_unit_0_register_file_0_n_145), .A(
      execution_unit_0_register_file_0_n_66_4));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r10_reg[3] (.Q(
      execution_unit_0_register_file_0_r10[3]), .QN(), .CK(
      execution_unit_0_register_file_0_n_141), .D(
      execution_unit_0_register_file_0_n_145), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_70 (.ZN(
      execution_unit_0_register_file_0_n_105_67), .A1(
      execution_unit_0_register_file_0_n_140), .A2(
      execution_unit_0_register_file_0_r10[3]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_59_7 (.ZN(
      execution_unit_0_register_file_0_n_59_4), .A1(
      execution_unit_0_register_file_0_n_59_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[3]), .B1(
      execution_unit_0_register_file_0_r9_wr), .B2(execution_unit_0_alu_out[3]));
  INV_X1_LVT execution_unit_0_register_file_0_i_59_8 (.ZN(
      execution_unit_0_register_file_0_n_126), .A(
      execution_unit_0_register_file_0_n_59_4));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r9_reg[3] (.Q(
      execution_unit_0_register_file_0_r9[3]), .QN(), .CK(
      execution_unit_0_register_file_0_n_122), .D(
      execution_unit_0_register_file_0_n_126), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_71 (.ZN(
      execution_unit_0_register_file_0_n_105_68), .A1(
      execution_unit_0_register_file_0_n_121), .A2(
      execution_unit_0_register_file_0_r9[3]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_105_72 (.ZN(
      execution_unit_0_register_file_0_n_105_69), .A1(
      execution_unit_0_register_file_0_n_105_65), .A2(
      execution_unit_0_register_file_0_n_105_66), .A3(
      execution_unit_0_register_file_0_n_105_67), .A4(
      execution_unit_0_register_file_0_n_105_68));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_52_7 (.ZN(
      execution_unit_0_register_file_0_n_52_4), .A1(
      execution_unit_0_register_file_0_n_52_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[3]), .B1(
      execution_unit_0_register_file_0_r8_wr), .B2(execution_unit_0_alu_out[3]));
  INV_X1_LVT execution_unit_0_register_file_0_i_52_8 (.ZN(
      execution_unit_0_register_file_0_n_107), .A(
      execution_unit_0_register_file_0_n_52_4));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r8_reg[3] (.Q(
      execution_unit_0_register_file_0_r8[3]), .QN(), .CK(
      execution_unit_0_register_file_0_n_103), .D(
      execution_unit_0_register_file_0_n_107), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_73 (.ZN(
      execution_unit_0_register_file_0_n_105_70), .A1(
      execution_unit_0_register_file_0_n_102), .A2(
      execution_unit_0_register_file_0_r8[3]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_45_7 (.ZN(
      execution_unit_0_register_file_0_n_45_4), .A1(
      execution_unit_0_register_file_0_n_45_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[3]), .B1(
      execution_unit_0_register_file_0_r7_wr), .B2(execution_unit_0_alu_out[3]));
  INV_X1_LVT execution_unit_0_register_file_0_i_45_8 (.ZN(
      execution_unit_0_register_file_0_n_88), .A(
      execution_unit_0_register_file_0_n_45_4));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r7_reg[3] (.Q(
      execution_unit_0_register_file_0_r7[3]), .QN(), .CK(
      execution_unit_0_register_file_0_n_84), .D(
      execution_unit_0_register_file_0_n_88), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_74 (.ZN(
      execution_unit_0_register_file_0_n_105_71), .A1(
      execution_unit_0_register_file_0_n_83), .A2(
      execution_unit_0_register_file_0_r7[3]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_38_7 (.ZN(
      execution_unit_0_register_file_0_n_38_4), .A1(
      execution_unit_0_register_file_0_n_38_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[3]), .B1(
      execution_unit_0_register_file_0_r6_wr), .B2(execution_unit_0_alu_out[3]));
  INV_X1_LVT execution_unit_0_register_file_0_i_38_8 (.ZN(
      execution_unit_0_register_file_0_n_69), .A(
      execution_unit_0_register_file_0_n_38_4));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r6_reg[3] (.Q(
      execution_unit_0_register_file_0_r6[3]), .QN(), .CK(
      execution_unit_0_register_file_0_n_65), .D(
      execution_unit_0_register_file_0_n_69), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_75 (.ZN(
      execution_unit_0_register_file_0_n_105_72), .A1(
      execution_unit_0_register_file_0_n_64), .A2(
      execution_unit_0_register_file_0_r6[3]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_31_7 (.ZN(
      execution_unit_0_register_file_0_n_31_4), .A1(
      execution_unit_0_register_file_0_n_31_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[3]), .B1(
      execution_unit_0_register_file_0_r5_wr), .B2(execution_unit_0_alu_out[3]));
  INV_X1_LVT execution_unit_0_register_file_0_i_31_8 (.ZN(
      execution_unit_0_register_file_0_n_50), .A(
      execution_unit_0_register_file_0_n_31_4));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r5_reg[3] (.Q(
      execution_unit_0_register_file_0_r5[3]), .QN(), .CK(
      execution_unit_0_register_file_0_n_46), .D(
      execution_unit_0_register_file_0_n_50), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_76 (.ZN(
      execution_unit_0_register_file_0_n_105_73), .A1(
      execution_unit_0_register_file_0_n_45), .A2(
      execution_unit_0_register_file_0_r5[3]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_105_77 (.ZN(
      execution_unit_0_register_file_0_n_105_74), .A1(
      execution_unit_0_register_file_0_n_105_70), .A2(
      execution_unit_0_register_file_0_n_105_71), .A3(
      execution_unit_0_register_file_0_n_105_72), .A4(
      execution_unit_0_register_file_0_n_105_73));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_87_7 (.ZN(
      execution_unit_0_register_file_0_n_87_4), .A1(
      execution_unit_0_register_file_0_n_87_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[3]), .B1(
      execution_unit_0_register_file_0_r13_wr), .B2(execution_unit_0_alu_out[3]));
  INV_X1_LVT execution_unit_0_register_file_0_i_87_8 (.ZN(
      execution_unit_0_register_file_0_n_202), .A(
      execution_unit_0_register_file_0_n_87_4));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r13_reg[3] (.Q(
      execution_unit_0_register_file_0_r13[3]), .QN(), .CK(
      execution_unit_0_register_file_0_n_198), .D(
      execution_unit_0_register_file_0_n_202), .RN(
      execution_unit_0_register_file_0_n_8));
  AND2_X1_LVT execution_unit_0_register_file_0_i_105_78 (.ZN(
      execution_unit_0_register_file_0_n_105_75), .A1(
      execution_unit_0_register_file_0_n_197), .A2(
      execution_unit_0_register_file_0_r13[3]));
  NOR4_X1_LVT execution_unit_0_register_file_0_i_105_79 (.ZN(
      execution_unit_0_register_file_0_n_105_76), .A1(
      execution_unit_0_register_file_0_n_105_64), .A2(
      execution_unit_0_register_file_0_n_105_69), .A3(
      execution_unit_0_register_file_0_n_105_74), .A4(
      execution_unit_0_register_file_0_n_105_75));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_80 (.ZN(
      execution_unit_0_register_file_0_n_105_77), .A1(
      execution_unit_0_register_file_0_n_254), .A2(pc[3]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_101_7 (.ZN(
      execution_unit_0_register_file_0_n_101_4), .A1(
      execution_unit_0_register_file_0_n_101_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[3]), .B1(
      execution_unit_0_register_file_0_r15_wr), .B2(execution_unit_0_alu_out[3]));
  INV_X1_LVT execution_unit_0_register_file_0_i_101_8 (.ZN(
      execution_unit_0_register_file_0_n_240), .A(
      execution_unit_0_register_file_0_n_101_4));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r15_reg[3] (.Q(
      execution_unit_0_register_file_0_r15[3]), .QN(), .CK(
      execution_unit_0_register_file_0_n_236), .D(
      execution_unit_0_register_file_0_n_240), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_81 (.ZN(
      execution_unit_0_register_file_0_n_105_78), .A1(
      execution_unit_0_register_file_0_n_235), .A2(
      execution_unit_0_register_file_0_r15[3]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_94_7 (.ZN(
      execution_unit_0_register_file_0_n_94_4), .A1(
      execution_unit_0_register_file_0_n_94_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[3]), .B1(
      execution_unit_0_register_file_0_r14_wr), .B2(execution_unit_0_alu_out[3]));
  INV_X1_LVT execution_unit_0_register_file_0_i_94_8 (.ZN(
      execution_unit_0_register_file_0_n_221), .A(
      execution_unit_0_register_file_0_n_94_4));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r14_reg[3] (.Q(
      execution_unit_0_register_file_0_r14[3]), .QN(), .CK(
      execution_unit_0_register_file_0_n_217), .D(
      execution_unit_0_register_file_0_n_221), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_82 (.ZN(
      execution_unit_0_register_file_0_n_105_79), .A1(
      execution_unit_0_register_file_0_n_216), .A2(
      execution_unit_0_register_file_0_r14[3]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_105_83 (.ZN(
      execution_unit_0_reg_src[3]), .A1(
      execution_unit_0_register_file_0_n_105_76), .A2(
      execution_unit_0_register_file_0_n_105_77), .A3(
      execution_unit_0_register_file_0_n_105_78), .A4(
      execution_unit_0_register_file_0_n_105_79));
  HA_X1_LVT execution_unit_0_register_file_0_i_22_3 (.CO(
      execution_unit_0_register_file_0_n_22_3), .S(
      execution_unit_0_register_file_0_reg_incr_val[3]), .A(
      execution_unit_0_reg_src[3]), .B(execution_unit_0_register_file_0_n_22_2));
  HA_X1_LVT execution_unit_0_register_file_0_i_22_4 (.CO(
      execution_unit_0_register_file_0_n_22_4), .S(
      execution_unit_0_register_file_0_reg_incr_val[4]), .A(
      execution_unit_0_reg_src[4]), .B(execution_unit_0_register_file_0_n_22_3));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_24_9 (.ZN(
      execution_unit_0_register_file_0_n_24_5), .A1(
      execution_unit_0_register_file_0_n_24_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[4]), .B1(
      execution_unit_0_register_file_0_r4_wr), .B2(execution_unit_0_alu_out[4]));
  INV_X1_LVT execution_unit_0_register_file_0_i_24_10 (.ZN(
      execution_unit_0_register_file_0_n_32), .A(
      execution_unit_0_register_file_0_n_24_5));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r4_reg[4] (.Q(
      execution_unit_0_register_file_0_r4[4]), .QN(), .CK(
      execution_unit_0_register_file_0_n_27), .D(
      execution_unit_0_register_file_0_n_32), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_84 (.ZN(
      execution_unit_0_register_file_0_n_105_80), .A1(
      execution_unit_0_register_file_0_n_24), .A2(
      execution_unit_0_register_file_0_r4[4]));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r3_reg[4] (.Q(
      execution_unit_0_register_file_0_r3[4]), .QN(), .CK(
      execution_unit_0_register_file_0_n_23), .D(execution_unit_0_alu_out[4]), 
      .RN(execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_85 (.ZN(
      execution_unit_0_register_file_0_n_105_81), .A1(
      execution_unit_0_register_file_0_n_22), .A2(
      execution_unit_0_register_file_0_r3[4]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_86 (.ZN(
      execution_unit_0_register_file_0_n_105_82), .A1(
      execution_unit_0_register_file_0_n_21), .A2(
      execution_unit_0_register_file_0_n_7));
  AOI222_X1_LVT execution_unit_0_register_file_0_i_109_6 (.ZN(
      execution_unit_0_register_file_0_n_109_3), .A1(
      execution_unit_0_register_file_0_r1_wr), .A2(execution_unit_0_alu_out[4]), 
      .B1(execution_unit_0_register_file_0_n_272), .B2(eu_mab[4]), .C1(
      execution_unit_0_register_file_0_n_271), .C2(
      execution_unit_0_register_file_0_n_258));
  INV_X1_LVT execution_unit_0_register_file_0_i_109_7 (.ZN(
      execution_unit_0_register_file_0_n_276), .A(
      execution_unit_0_register_file_0_n_109_3));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r1_reg[4] (.Q(
      execution_unit_0_register_file_0_r1[4]), .QN(), .CK(
      execution_unit_0_register_file_0_n_270), .D(
      execution_unit_0_register_file_0_n_276), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_87 (.ZN(
      execution_unit_0_register_file_0_n_105_83), .A1(
      execution_unit_0_register_file_0_inst_src_in), .A2(
      execution_unit_0_register_file_0_r1[4]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_105_88 (.ZN(
      execution_unit_0_register_file_0_n_105_84), .A1(
      execution_unit_0_register_file_0_n_105_80), .A2(
      execution_unit_0_register_file_0_n_105_81), .A3(
      execution_unit_0_register_file_0_n_105_82), .A4(
      execution_unit_0_register_file_0_n_105_83));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_80_9 (.ZN(
      execution_unit_0_register_file_0_n_80_5), .A1(
      execution_unit_0_register_file_0_n_80_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[4]), .B1(
      execution_unit_0_register_file_0_r12_wr), .B2(execution_unit_0_alu_out[4]));
  INV_X1_LVT execution_unit_0_register_file_0_i_80_10 (.ZN(
      execution_unit_0_register_file_0_n_184), .A(
      execution_unit_0_register_file_0_n_80_5));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r12_reg[4] (.Q(
      execution_unit_0_register_file_0_r12[4]), .QN(), .CK(
      execution_unit_0_register_file_0_n_179), .D(
      execution_unit_0_register_file_0_n_184), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_89 (.ZN(
      execution_unit_0_register_file_0_n_105_85), .A1(
      execution_unit_0_register_file_0_n_178), .A2(
      execution_unit_0_register_file_0_r12[4]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_73_9 (.ZN(
      execution_unit_0_register_file_0_n_73_5), .A1(
      execution_unit_0_register_file_0_n_73_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[4]), .B1(
      execution_unit_0_register_file_0_r11_wr), .B2(execution_unit_0_alu_out[4]));
  INV_X1_LVT execution_unit_0_register_file_0_i_73_10 (.ZN(
      execution_unit_0_register_file_0_n_165), .A(
      execution_unit_0_register_file_0_n_73_5));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r11_reg[4] (.Q(
      execution_unit_0_register_file_0_r11[4]), .QN(), .CK(
      execution_unit_0_register_file_0_n_160), .D(
      execution_unit_0_register_file_0_n_165), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_90 (.ZN(
      execution_unit_0_register_file_0_n_105_86), .A1(
      execution_unit_0_register_file_0_n_159), .A2(
      execution_unit_0_register_file_0_r11[4]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_66_9 (.ZN(
      execution_unit_0_register_file_0_n_66_5), .A1(
      execution_unit_0_register_file_0_n_66_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[4]), .B1(
      execution_unit_0_register_file_0_r10_wr), .B2(execution_unit_0_alu_out[4]));
  INV_X1_LVT execution_unit_0_register_file_0_i_66_10 (.ZN(
      execution_unit_0_register_file_0_n_146), .A(
      execution_unit_0_register_file_0_n_66_5));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r10_reg[4] (.Q(
      execution_unit_0_register_file_0_r10[4]), .QN(), .CK(
      execution_unit_0_register_file_0_n_141), .D(
      execution_unit_0_register_file_0_n_146), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_91 (.ZN(
      execution_unit_0_register_file_0_n_105_87), .A1(
      execution_unit_0_register_file_0_n_140), .A2(
      execution_unit_0_register_file_0_r10[4]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_59_9 (.ZN(
      execution_unit_0_register_file_0_n_59_5), .A1(
      execution_unit_0_register_file_0_n_59_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[4]), .B1(
      execution_unit_0_register_file_0_r9_wr), .B2(execution_unit_0_alu_out[4]));
  INV_X1_LVT execution_unit_0_register_file_0_i_59_10 (.ZN(
      execution_unit_0_register_file_0_n_127), .A(
      execution_unit_0_register_file_0_n_59_5));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r9_reg[4] (.Q(
      execution_unit_0_register_file_0_r9[4]), .QN(), .CK(
      execution_unit_0_register_file_0_n_122), .D(
      execution_unit_0_register_file_0_n_127), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_92 (.ZN(
      execution_unit_0_register_file_0_n_105_88), .A1(
      execution_unit_0_register_file_0_n_121), .A2(
      execution_unit_0_register_file_0_r9[4]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_105_93 (.ZN(
      execution_unit_0_register_file_0_n_105_89), .A1(
      execution_unit_0_register_file_0_n_105_85), .A2(
      execution_unit_0_register_file_0_n_105_86), .A3(
      execution_unit_0_register_file_0_n_105_87), .A4(
      execution_unit_0_register_file_0_n_105_88));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_52_9 (.ZN(
      execution_unit_0_register_file_0_n_52_5), .A1(
      execution_unit_0_register_file_0_n_52_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[4]), .B1(
      execution_unit_0_register_file_0_r8_wr), .B2(execution_unit_0_alu_out[4]));
  INV_X1_LVT execution_unit_0_register_file_0_i_52_10 (.ZN(
      execution_unit_0_register_file_0_n_108), .A(
      execution_unit_0_register_file_0_n_52_5));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r8_reg[4] (.Q(
      execution_unit_0_register_file_0_r8[4]), .QN(), .CK(
      execution_unit_0_register_file_0_n_103), .D(
      execution_unit_0_register_file_0_n_108), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_94 (.ZN(
      execution_unit_0_register_file_0_n_105_90), .A1(
      execution_unit_0_register_file_0_n_102), .A2(
      execution_unit_0_register_file_0_r8[4]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_45_9 (.ZN(
      execution_unit_0_register_file_0_n_45_5), .A1(
      execution_unit_0_register_file_0_n_45_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[4]), .B1(
      execution_unit_0_register_file_0_r7_wr), .B2(execution_unit_0_alu_out[4]));
  INV_X1_LVT execution_unit_0_register_file_0_i_45_10 (.ZN(
      execution_unit_0_register_file_0_n_89), .A(
      execution_unit_0_register_file_0_n_45_5));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r7_reg[4] (.Q(
      execution_unit_0_register_file_0_r7[4]), .QN(), .CK(
      execution_unit_0_register_file_0_n_84), .D(
      execution_unit_0_register_file_0_n_89), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_95 (.ZN(
      execution_unit_0_register_file_0_n_105_91), .A1(
      execution_unit_0_register_file_0_n_83), .A2(
      execution_unit_0_register_file_0_r7[4]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_38_9 (.ZN(
      execution_unit_0_register_file_0_n_38_5), .A1(
      execution_unit_0_register_file_0_n_38_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[4]), .B1(
      execution_unit_0_register_file_0_r6_wr), .B2(execution_unit_0_alu_out[4]));
  INV_X1_LVT execution_unit_0_register_file_0_i_38_10 (.ZN(
      execution_unit_0_register_file_0_n_70), .A(
      execution_unit_0_register_file_0_n_38_5));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r6_reg[4] (.Q(
      execution_unit_0_register_file_0_r6[4]), .QN(), .CK(
      execution_unit_0_register_file_0_n_65), .D(
      execution_unit_0_register_file_0_n_70), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_96 (.ZN(
      execution_unit_0_register_file_0_n_105_92), .A1(
      execution_unit_0_register_file_0_n_64), .A2(
      execution_unit_0_register_file_0_r6[4]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_31_9 (.ZN(
      execution_unit_0_register_file_0_n_31_5), .A1(
      execution_unit_0_register_file_0_n_31_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[4]), .B1(
      execution_unit_0_register_file_0_r5_wr), .B2(execution_unit_0_alu_out[4]));
  INV_X1_LVT execution_unit_0_register_file_0_i_31_10 (.ZN(
      execution_unit_0_register_file_0_n_51), .A(
      execution_unit_0_register_file_0_n_31_5));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r5_reg[4] (.Q(
      execution_unit_0_register_file_0_r5[4]), .QN(), .CK(
      execution_unit_0_register_file_0_n_46), .D(
      execution_unit_0_register_file_0_n_51), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_97 (.ZN(
      execution_unit_0_register_file_0_n_105_93), .A1(
      execution_unit_0_register_file_0_n_45), .A2(
      execution_unit_0_register_file_0_r5[4]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_105_98 (.ZN(
      execution_unit_0_register_file_0_n_105_94), .A1(
      execution_unit_0_register_file_0_n_105_90), .A2(
      execution_unit_0_register_file_0_n_105_91), .A3(
      execution_unit_0_register_file_0_n_105_92), .A4(
      execution_unit_0_register_file_0_n_105_93));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_87_9 (.ZN(
      execution_unit_0_register_file_0_n_87_5), .A1(
      execution_unit_0_register_file_0_n_87_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[4]), .B1(
      execution_unit_0_register_file_0_r13_wr), .B2(execution_unit_0_alu_out[4]));
  INV_X1_LVT execution_unit_0_register_file_0_i_87_10 (.ZN(
      execution_unit_0_register_file_0_n_203), .A(
      execution_unit_0_register_file_0_n_87_5));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r13_reg[4] (.Q(
      execution_unit_0_register_file_0_r13[4]), .QN(), .CK(
      execution_unit_0_register_file_0_n_198), .D(
      execution_unit_0_register_file_0_n_203), .RN(
      execution_unit_0_register_file_0_n_8));
  AND2_X1_LVT execution_unit_0_register_file_0_i_105_99 (.ZN(
      execution_unit_0_register_file_0_n_105_95), .A1(
      execution_unit_0_register_file_0_n_197), .A2(
      execution_unit_0_register_file_0_r13[4]));
  NOR4_X1_LVT execution_unit_0_register_file_0_i_105_100 (.ZN(
      execution_unit_0_register_file_0_n_105_96), .A1(
      execution_unit_0_register_file_0_n_105_84), .A2(
      execution_unit_0_register_file_0_n_105_89), .A3(
      execution_unit_0_register_file_0_n_105_94), .A4(
      execution_unit_0_register_file_0_n_105_95));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_101 (.ZN(
      execution_unit_0_register_file_0_n_105_97), .A1(
      execution_unit_0_register_file_0_n_254), .A2(pc[4]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_101_9 (.ZN(
      execution_unit_0_register_file_0_n_101_5), .A1(
      execution_unit_0_register_file_0_n_101_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[4]), .B1(
      execution_unit_0_register_file_0_r15_wr), .B2(execution_unit_0_alu_out[4]));
  INV_X1_LVT execution_unit_0_register_file_0_i_101_10 (.ZN(
      execution_unit_0_register_file_0_n_241), .A(
      execution_unit_0_register_file_0_n_101_5));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r15_reg[4] (.Q(
      execution_unit_0_register_file_0_r15[4]), .QN(), .CK(
      execution_unit_0_register_file_0_n_236), .D(
      execution_unit_0_register_file_0_n_241), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_102 (.ZN(
      execution_unit_0_register_file_0_n_105_98), .A1(
      execution_unit_0_register_file_0_n_235), .A2(
      execution_unit_0_register_file_0_r15[4]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_94_9 (.ZN(
      execution_unit_0_register_file_0_n_94_5), .A1(
      execution_unit_0_register_file_0_n_94_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[4]), .B1(
      execution_unit_0_register_file_0_r14_wr), .B2(execution_unit_0_alu_out[4]));
  INV_X1_LVT execution_unit_0_register_file_0_i_94_10 (.ZN(
      execution_unit_0_register_file_0_n_222), .A(
      execution_unit_0_register_file_0_n_94_5));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r14_reg[4] (.Q(
      execution_unit_0_register_file_0_r14[4]), .QN(), .CK(
      execution_unit_0_register_file_0_n_217), .D(
      execution_unit_0_register_file_0_n_222), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_103 (.ZN(
      execution_unit_0_register_file_0_n_105_99), .A1(
      execution_unit_0_register_file_0_n_216), .A2(
      execution_unit_0_register_file_0_r14[4]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_105_104 (.ZN(
      execution_unit_0_reg_src[4]), .A1(
      execution_unit_0_register_file_0_n_105_96), .A2(
      execution_unit_0_register_file_0_n_105_97), .A3(
      execution_unit_0_register_file_0_n_105_98), .A4(
      execution_unit_0_register_file_0_n_105_99));
  HA_X1_LVT execution_unit_0_register_file_0_i_106_3 (.CO(
      execution_unit_0_register_file_0_n_106_2), .S(
      execution_unit_0_register_file_0_n_258), .A(execution_unit_0_reg_src[4]), 
      .B(execution_unit_0_register_file_0_n_106_1));
  HA_X1_LVT execution_unit_0_register_file_0_i_106_4 (.CO(
      execution_unit_0_register_file_0_n_106_3), .S(
      execution_unit_0_register_file_0_n_259), .A(execution_unit_0_reg_src[5]), 
      .B(execution_unit_0_register_file_0_n_106_2));
  AOI222_X1_LVT execution_unit_0_register_file_0_i_109_8 (.ZN(
      execution_unit_0_register_file_0_n_109_4), .A1(
      execution_unit_0_register_file_0_r1_wr), .A2(execution_unit_0_alu_out[5]), 
      .B1(execution_unit_0_register_file_0_n_272), .B2(eu_mab[5]), .C1(
      execution_unit_0_register_file_0_n_271), .C2(
      execution_unit_0_register_file_0_n_259));
  INV_X1_LVT execution_unit_0_register_file_0_i_109_9 (.ZN(
      execution_unit_0_register_file_0_n_277), .A(
      execution_unit_0_register_file_0_n_109_4));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r1_reg[5] (.Q(
      execution_unit_0_register_file_0_r1[5]), .QN(), .CK(
      execution_unit_0_register_file_0_n_270), .D(
      execution_unit_0_register_file_0_n_277), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_108 (.ZN(
      execution_unit_0_register_file_0_n_105_103), .A1(
      execution_unit_0_register_file_0_inst_src_in), .A2(
      execution_unit_0_register_file_0_r1[5]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_105_109 (.ZN(
      execution_unit_0_register_file_0_n_105_104), .A1(
      execution_unit_0_register_file_0_n_105_100), .A2(
      execution_unit_0_register_file_0_n_105_101), .A3(
      execution_unit_0_register_file_0_n_105_102), .A4(
      execution_unit_0_register_file_0_n_105_103));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_80_11 (.ZN(
      execution_unit_0_register_file_0_n_80_6), .A1(
      execution_unit_0_register_file_0_n_80_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[5]), .B1(
      execution_unit_0_register_file_0_r12_wr), .B2(execution_unit_0_alu_out[5]));
  INV_X1_LVT execution_unit_0_register_file_0_i_80_12 (.ZN(
      execution_unit_0_register_file_0_n_185), .A(
      execution_unit_0_register_file_0_n_80_6));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r12_reg[5] (.Q(
      execution_unit_0_register_file_0_r12[5]), .QN(), .CK(
      execution_unit_0_register_file_0_n_179), .D(
      execution_unit_0_register_file_0_n_185), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_110 (.ZN(
      execution_unit_0_register_file_0_n_105_105), .A1(
      execution_unit_0_register_file_0_n_178), .A2(
      execution_unit_0_register_file_0_r12[5]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_73_11 (.ZN(
      execution_unit_0_register_file_0_n_73_6), .A1(
      execution_unit_0_register_file_0_n_73_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[5]), .B1(
      execution_unit_0_register_file_0_r11_wr), .B2(execution_unit_0_alu_out[5]));
  INV_X1_LVT execution_unit_0_register_file_0_i_73_12 (.ZN(
      execution_unit_0_register_file_0_n_166), .A(
      execution_unit_0_register_file_0_n_73_6));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r11_reg[5] (.Q(
      execution_unit_0_register_file_0_r11[5]), .QN(), .CK(
      execution_unit_0_register_file_0_n_160), .D(
      execution_unit_0_register_file_0_n_166), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_111 (.ZN(
      execution_unit_0_register_file_0_n_105_106), .A1(
      execution_unit_0_register_file_0_n_159), .A2(
      execution_unit_0_register_file_0_r11[5]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_66_11 (.ZN(
      execution_unit_0_register_file_0_n_66_6), .A1(
      execution_unit_0_register_file_0_n_66_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[5]), .B1(
      execution_unit_0_register_file_0_r10_wr), .B2(execution_unit_0_alu_out[5]));
  INV_X1_LVT execution_unit_0_register_file_0_i_66_12 (.ZN(
      execution_unit_0_register_file_0_n_147), .A(
      execution_unit_0_register_file_0_n_66_6));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r10_reg[5] (.Q(
      execution_unit_0_register_file_0_r10[5]), .QN(), .CK(
      execution_unit_0_register_file_0_n_141), .D(
      execution_unit_0_register_file_0_n_147), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_112 (.ZN(
      execution_unit_0_register_file_0_n_105_107), .A1(
      execution_unit_0_register_file_0_n_140), .A2(
      execution_unit_0_register_file_0_r10[5]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_59_11 (.ZN(
      execution_unit_0_register_file_0_n_59_6), .A1(
      execution_unit_0_register_file_0_n_59_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[5]), .B1(
      execution_unit_0_register_file_0_r9_wr), .B2(execution_unit_0_alu_out[5]));
  INV_X1_LVT execution_unit_0_register_file_0_i_59_12 (.ZN(
      execution_unit_0_register_file_0_n_128), .A(
      execution_unit_0_register_file_0_n_59_6));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r9_reg[5] (.Q(
      execution_unit_0_register_file_0_r9[5]), .QN(), .CK(
      execution_unit_0_register_file_0_n_122), .D(
      execution_unit_0_register_file_0_n_128), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_113 (.ZN(
      execution_unit_0_register_file_0_n_105_108), .A1(
      execution_unit_0_register_file_0_n_121), .A2(
      execution_unit_0_register_file_0_r9[5]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_105_114 (.ZN(
      execution_unit_0_register_file_0_n_105_109), .A1(
      execution_unit_0_register_file_0_n_105_105), .A2(
      execution_unit_0_register_file_0_n_105_106), .A3(
      execution_unit_0_register_file_0_n_105_107), .A4(
      execution_unit_0_register_file_0_n_105_108));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_52_11 (.ZN(
      execution_unit_0_register_file_0_n_52_6), .A1(
      execution_unit_0_register_file_0_n_52_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[5]), .B1(
      execution_unit_0_register_file_0_r8_wr), .B2(execution_unit_0_alu_out[5]));
  INV_X1_LVT execution_unit_0_register_file_0_i_52_12 (.ZN(
      execution_unit_0_register_file_0_n_109), .A(
      execution_unit_0_register_file_0_n_52_6));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r8_reg[5] (.Q(
      execution_unit_0_register_file_0_r8[5]), .QN(), .CK(
      execution_unit_0_register_file_0_n_103), .D(
      execution_unit_0_register_file_0_n_109), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_115 (.ZN(
      execution_unit_0_register_file_0_n_105_110), .A1(
      execution_unit_0_register_file_0_n_102), .A2(
      execution_unit_0_register_file_0_r8[5]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_45_11 (.ZN(
      execution_unit_0_register_file_0_n_45_6), .A1(
      execution_unit_0_register_file_0_n_45_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[5]), .B1(
      execution_unit_0_register_file_0_r7_wr), .B2(execution_unit_0_alu_out[5]));
  INV_X1_LVT execution_unit_0_register_file_0_i_45_12 (.ZN(
      execution_unit_0_register_file_0_n_90), .A(
      execution_unit_0_register_file_0_n_45_6));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r7_reg[5] (.Q(
      execution_unit_0_register_file_0_r7[5]), .QN(), .CK(
      execution_unit_0_register_file_0_n_84), .D(
      execution_unit_0_register_file_0_n_90), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_116 (.ZN(
      execution_unit_0_register_file_0_n_105_111), .A1(
      execution_unit_0_register_file_0_n_83), .A2(
      execution_unit_0_register_file_0_r7[5]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_38_11 (.ZN(
      execution_unit_0_register_file_0_n_38_6), .A1(
      execution_unit_0_register_file_0_n_38_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[5]), .B1(
      execution_unit_0_register_file_0_r6_wr), .B2(execution_unit_0_alu_out[5]));
  INV_X1_LVT execution_unit_0_register_file_0_i_38_12 (.ZN(
      execution_unit_0_register_file_0_n_71), .A(
      execution_unit_0_register_file_0_n_38_6));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r6_reg[5] (.Q(
      execution_unit_0_register_file_0_r6[5]), .QN(), .CK(
      execution_unit_0_register_file_0_n_65), .D(
      execution_unit_0_register_file_0_n_71), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_117 (.ZN(
      execution_unit_0_register_file_0_n_105_112), .A1(
      execution_unit_0_register_file_0_n_64), .A2(
      execution_unit_0_register_file_0_r6[5]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_31_11 (.ZN(
      execution_unit_0_register_file_0_n_31_6), .A1(
      execution_unit_0_register_file_0_n_31_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[5]), .B1(
      execution_unit_0_register_file_0_r5_wr), .B2(execution_unit_0_alu_out[5]));
  INV_X1_LVT execution_unit_0_register_file_0_i_31_12 (.ZN(
      execution_unit_0_register_file_0_n_52), .A(
      execution_unit_0_register_file_0_n_31_6));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r5_reg[5] (.Q(
      execution_unit_0_register_file_0_r5[5]), .QN(), .CK(
      execution_unit_0_register_file_0_n_46), .D(
      execution_unit_0_register_file_0_n_52), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_118 (.ZN(
      execution_unit_0_register_file_0_n_105_113), .A1(
      execution_unit_0_register_file_0_n_45), .A2(
      execution_unit_0_register_file_0_r5[5]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_105_119 (.ZN(
      execution_unit_0_register_file_0_n_105_114), .A1(
      execution_unit_0_register_file_0_n_105_110), .A2(
      execution_unit_0_register_file_0_n_105_111), .A3(
      execution_unit_0_register_file_0_n_105_112), .A4(
      execution_unit_0_register_file_0_n_105_113));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_87_11 (.ZN(
      execution_unit_0_register_file_0_n_87_6), .A1(
      execution_unit_0_register_file_0_n_87_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[5]), .B1(
      execution_unit_0_register_file_0_r13_wr), .B2(execution_unit_0_alu_out[5]));
  INV_X1_LVT execution_unit_0_register_file_0_i_87_12 (.ZN(
      execution_unit_0_register_file_0_n_204), .A(
      execution_unit_0_register_file_0_n_87_6));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r13_reg[5] (.Q(
      execution_unit_0_register_file_0_r13[5]), .QN(), .CK(
      execution_unit_0_register_file_0_n_198), .D(
      execution_unit_0_register_file_0_n_204), .RN(
      execution_unit_0_register_file_0_n_8));
  AND2_X1_LVT execution_unit_0_register_file_0_i_105_120 (.ZN(
      execution_unit_0_register_file_0_n_105_115), .A1(
      execution_unit_0_register_file_0_n_197), .A2(
      execution_unit_0_register_file_0_r13[5]));
  NOR4_X1_LVT execution_unit_0_register_file_0_i_105_121 (.ZN(
      execution_unit_0_register_file_0_n_105_116), .A1(
      execution_unit_0_register_file_0_n_105_104), .A2(
      execution_unit_0_register_file_0_n_105_109), .A3(
      execution_unit_0_register_file_0_n_105_114), .A4(
      execution_unit_0_register_file_0_n_105_115));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_122 (.ZN(
      execution_unit_0_register_file_0_n_105_117), .A1(
      execution_unit_0_register_file_0_n_254), .A2(pc[5]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_101_11 (.ZN(
      execution_unit_0_register_file_0_n_101_6), .A1(
      execution_unit_0_register_file_0_n_101_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[5]), .B1(
      execution_unit_0_register_file_0_r15_wr), .B2(execution_unit_0_alu_out[5]));
  INV_X1_LVT execution_unit_0_register_file_0_i_101_12 (.ZN(
      execution_unit_0_register_file_0_n_242), .A(
      execution_unit_0_register_file_0_n_101_6));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r15_reg[5] (.Q(
      execution_unit_0_register_file_0_r15[5]), .QN(), .CK(
      execution_unit_0_register_file_0_n_236), .D(
      execution_unit_0_register_file_0_n_242), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_123 (.ZN(
      execution_unit_0_register_file_0_n_105_118), .A1(
      execution_unit_0_register_file_0_n_235), .A2(
      execution_unit_0_register_file_0_r15[5]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_94_11 (.ZN(
      execution_unit_0_register_file_0_n_94_6), .A1(
      execution_unit_0_register_file_0_n_94_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[5]), .B1(
      execution_unit_0_register_file_0_r14_wr), .B2(execution_unit_0_alu_out[5]));
  INV_X1_LVT execution_unit_0_register_file_0_i_94_12 (.ZN(
      execution_unit_0_register_file_0_n_223), .A(
      execution_unit_0_register_file_0_n_94_6));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r14_reg[5] (.Q(
      execution_unit_0_register_file_0_r14[5]), .QN(), .CK(
      execution_unit_0_register_file_0_n_217), .D(
      execution_unit_0_register_file_0_n_223), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_124 (.ZN(
      execution_unit_0_register_file_0_n_105_119), .A1(
      execution_unit_0_register_file_0_n_216), .A2(
      execution_unit_0_register_file_0_r14[5]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_105_125 (.ZN(
      execution_unit_0_reg_src[5]), .A1(
      execution_unit_0_register_file_0_n_105_116), .A2(
      execution_unit_0_register_file_0_n_105_117), .A3(
      execution_unit_0_register_file_0_n_105_118), .A4(
      execution_unit_0_register_file_0_n_105_119));
  HA_X1_LVT execution_unit_0_register_file_0_i_22_5 (.CO(
      execution_unit_0_register_file_0_n_22_5), .S(
      execution_unit_0_register_file_0_reg_incr_val[5]), .A(
      execution_unit_0_reg_src[5]), .B(execution_unit_0_register_file_0_n_22_4));
  HA_X1_LVT execution_unit_0_register_file_0_i_22_6 (.CO(
      execution_unit_0_register_file_0_n_22_6), .S(
      execution_unit_0_register_file_0_reg_incr_val[6]), .A(
      execution_unit_0_reg_src[6]), .B(execution_unit_0_register_file_0_n_22_5));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_24_13 (.ZN(
      execution_unit_0_register_file_0_n_24_7), .A1(
      execution_unit_0_register_file_0_n_24_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[6]), .B1(
      execution_unit_0_register_file_0_r4_wr), .B2(execution_unit_0_alu_out[6]));
  INV_X1_LVT execution_unit_0_register_file_0_i_24_14 (.ZN(
      execution_unit_0_register_file_0_n_34), .A(
      execution_unit_0_register_file_0_n_24_7));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r4_reg[6] (.Q(
      execution_unit_0_register_file_0_r4[6]), .QN(), .CK(
      execution_unit_0_register_file_0_n_27), .D(
      execution_unit_0_register_file_0_n_34), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_126 (.ZN(
      execution_unit_0_register_file_0_n_105_120), .A1(
      execution_unit_0_register_file_0_n_24), .A2(
      execution_unit_0_register_file_0_r4[6]));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r3_reg[6] (.Q(
      execution_unit_0_register_file_0_r3[6]), .QN(), .CK(
      execution_unit_0_register_file_0_n_23), .D(execution_unit_0_alu_out[6]), 
      .RN(execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_127 (.ZN(
      execution_unit_0_register_file_0_n_105_121), .A1(
      execution_unit_0_register_file_0_n_22), .A2(
      execution_unit_0_register_file_0_r3[6]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_2_5 (.ZN(
      execution_unit_0_register_file_0_n_2_3), .A1(
      execution_unit_0_register_file_0_n_2_0), .A2(scg0), .B1(
      execution_unit_0_register_file_0_r2_wr), .B2(execution_unit_0_alu_out[6]));
  INV_X1_LVT execution_unit_0_register_file_0_i_2_6 (.ZN(
      execution_unit_0_register_file_0_r2_nxt[3]), .A(
      execution_unit_0_register_file_0_n_2_3));
  AND2_X1_LVT execution_unit_0_register_file_0_i_6_6 (.ZN(
      execution_unit_0_register_file_0_n_18), .A1(
      execution_unit_0_register_file_0_n_6_0), .A2(
      execution_unit_0_register_file_0_r2_nxt[3]));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r2_reg[6] (.Q(scg0), .QN(), .CK(
      cpu_mclk), .D(execution_unit_0_register_file_0_n_18), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_128 (.ZN(
      execution_unit_0_register_file_0_n_105_122), .A1(
      execution_unit_0_register_file_0_n_21), .A2(scg0));
  AOI222_X1_LVT execution_unit_0_register_file_0_i_109_10 (.ZN(
      execution_unit_0_register_file_0_n_109_5), .A1(
      execution_unit_0_register_file_0_r1_wr), .A2(execution_unit_0_alu_out[6]), 
      .B1(execution_unit_0_register_file_0_n_272), .B2(eu_mab[6]), .C1(
      execution_unit_0_register_file_0_n_271), .C2(
      execution_unit_0_register_file_0_n_260));
  INV_X1_LVT execution_unit_0_register_file_0_i_109_11 (.ZN(
      execution_unit_0_register_file_0_n_278), .A(
      execution_unit_0_register_file_0_n_109_5));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r1_reg[6] (.Q(
      execution_unit_0_register_file_0_r1[6]), .QN(), .CK(
      execution_unit_0_register_file_0_n_270), .D(
      execution_unit_0_register_file_0_n_278), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_129 (.ZN(
      execution_unit_0_register_file_0_n_105_123), .A1(
      execution_unit_0_register_file_0_inst_src_in), .A2(
      execution_unit_0_register_file_0_r1[6]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_105_130 (.ZN(
      execution_unit_0_register_file_0_n_105_124), .A1(
      execution_unit_0_register_file_0_n_105_120), .A2(
      execution_unit_0_register_file_0_n_105_121), .A3(
      execution_unit_0_register_file_0_n_105_122), .A4(
      execution_unit_0_register_file_0_n_105_123));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_80_13 (.ZN(
      execution_unit_0_register_file_0_n_80_7), .A1(
      execution_unit_0_register_file_0_n_80_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[6]), .B1(
      execution_unit_0_register_file_0_r12_wr), .B2(execution_unit_0_alu_out[6]));
  INV_X1_LVT execution_unit_0_register_file_0_i_80_14 (.ZN(
      execution_unit_0_register_file_0_n_186), .A(
      execution_unit_0_register_file_0_n_80_7));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r12_reg[6] (.Q(
      execution_unit_0_register_file_0_r12[6]), .QN(), .CK(
      execution_unit_0_register_file_0_n_179), .D(
      execution_unit_0_register_file_0_n_186), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_131 (.ZN(
      execution_unit_0_register_file_0_n_105_125), .A1(
      execution_unit_0_register_file_0_n_178), .A2(
      execution_unit_0_register_file_0_r12[6]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_73_13 (.ZN(
      execution_unit_0_register_file_0_n_73_7), .A1(
      execution_unit_0_register_file_0_n_73_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[6]), .B1(
      execution_unit_0_register_file_0_r11_wr), .B2(execution_unit_0_alu_out[6]));
  INV_X1_LVT execution_unit_0_register_file_0_i_73_14 (.ZN(
      execution_unit_0_register_file_0_n_167), .A(
      execution_unit_0_register_file_0_n_73_7));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r11_reg[6] (.Q(
      execution_unit_0_register_file_0_r11[6]), .QN(), .CK(
      execution_unit_0_register_file_0_n_160), .D(
      execution_unit_0_register_file_0_n_167), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_132 (.ZN(
      execution_unit_0_register_file_0_n_105_126), .A1(
      execution_unit_0_register_file_0_n_159), .A2(
      execution_unit_0_register_file_0_r11[6]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_66_13 (.ZN(
      execution_unit_0_register_file_0_n_66_7), .A1(
      execution_unit_0_register_file_0_n_66_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[6]), .B1(
      execution_unit_0_register_file_0_r10_wr), .B2(execution_unit_0_alu_out[6]));
  INV_X1_LVT execution_unit_0_register_file_0_i_66_14 (.ZN(
      execution_unit_0_register_file_0_n_148), .A(
      execution_unit_0_register_file_0_n_66_7));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r10_reg[6] (.Q(
      execution_unit_0_register_file_0_r10[6]), .QN(), .CK(
      execution_unit_0_register_file_0_n_141), .D(
      execution_unit_0_register_file_0_n_148), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_133 (.ZN(
      execution_unit_0_register_file_0_n_105_127), .A1(
      execution_unit_0_register_file_0_n_140), .A2(
      execution_unit_0_register_file_0_r10[6]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_59_13 (.ZN(
      execution_unit_0_register_file_0_n_59_7), .A1(
      execution_unit_0_register_file_0_n_59_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[6]), .B1(
      execution_unit_0_register_file_0_r9_wr), .B2(execution_unit_0_alu_out[6]));
  INV_X1_LVT execution_unit_0_register_file_0_i_59_14 (.ZN(
      execution_unit_0_register_file_0_n_129), .A(
      execution_unit_0_register_file_0_n_59_7));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r9_reg[6] (.Q(
      execution_unit_0_register_file_0_r9[6]), .QN(), .CK(
      execution_unit_0_register_file_0_n_122), .D(
      execution_unit_0_register_file_0_n_129), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_134 (.ZN(
      execution_unit_0_register_file_0_n_105_128), .A1(
      execution_unit_0_register_file_0_n_121), .A2(
      execution_unit_0_register_file_0_r9[6]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_105_135 (.ZN(
      execution_unit_0_register_file_0_n_105_129), .A1(
      execution_unit_0_register_file_0_n_105_125), .A2(
      execution_unit_0_register_file_0_n_105_126), .A3(
      execution_unit_0_register_file_0_n_105_127), .A4(
      execution_unit_0_register_file_0_n_105_128));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_52_13 (.ZN(
      execution_unit_0_register_file_0_n_52_7), .A1(
      execution_unit_0_register_file_0_n_52_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[6]), .B1(
      execution_unit_0_register_file_0_r8_wr), .B2(execution_unit_0_alu_out[6]));
  INV_X1_LVT execution_unit_0_register_file_0_i_52_14 (.ZN(
      execution_unit_0_register_file_0_n_110), .A(
      execution_unit_0_register_file_0_n_52_7));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r8_reg[6] (.Q(
      execution_unit_0_register_file_0_r8[6]), .QN(), .CK(
      execution_unit_0_register_file_0_n_103), .D(
      execution_unit_0_register_file_0_n_110), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_136 (.ZN(
      execution_unit_0_register_file_0_n_105_130), .A1(
      execution_unit_0_register_file_0_n_102), .A2(
      execution_unit_0_register_file_0_r8[6]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_45_13 (.ZN(
      execution_unit_0_register_file_0_n_45_7), .A1(
      execution_unit_0_register_file_0_n_45_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[6]), .B1(
      execution_unit_0_register_file_0_r7_wr), .B2(execution_unit_0_alu_out[6]));
  INV_X1_LVT execution_unit_0_register_file_0_i_45_14 (.ZN(
      execution_unit_0_register_file_0_n_91), .A(
      execution_unit_0_register_file_0_n_45_7));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r7_reg[6] (.Q(
      execution_unit_0_register_file_0_r7[6]), .QN(), .CK(
      execution_unit_0_register_file_0_n_84), .D(
      execution_unit_0_register_file_0_n_91), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_137 (.ZN(
      execution_unit_0_register_file_0_n_105_131), .A1(
      execution_unit_0_register_file_0_n_83), .A2(
      execution_unit_0_register_file_0_r7[6]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_38_13 (.ZN(
      execution_unit_0_register_file_0_n_38_7), .A1(
      execution_unit_0_register_file_0_n_38_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[6]), .B1(
      execution_unit_0_register_file_0_r6_wr), .B2(execution_unit_0_alu_out[6]));
  INV_X1_LVT execution_unit_0_register_file_0_i_38_14 (.ZN(
      execution_unit_0_register_file_0_n_72), .A(
      execution_unit_0_register_file_0_n_38_7));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r6_reg[6] (.Q(
      execution_unit_0_register_file_0_r6[6]), .QN(), .CK(
      execution_unit_0_register_file_0_n_65), .D(
      execution_unit_0_register_file_0_n_72), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_138 (.ZN(
      execution_unit_0_register_file_0_n_105_132), .A1(
      execution_unit_0_register_file_0_n_64), .A2(
      execution_unit_0_register_file_0_r6[6]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_31_13 (.ZN(
      execution_unit_0_register_file_0_n_31_7), .A1(
      execution_unit_0_register_file_0_n_31_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[6]), .B1(
      execution_unit_0_register_file_0_r5_wr), .B2(execution_unit_0_alu_out[6]));
  INV_X1_LVT execution_unit_0_register_file_0_i_31_14 (.ZN(
      execution_unit_0_register_file_0_n_53), .A(
      execution_unit_0_register_file_0_n_31_7));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r5_reg[6] (.Q(
      execution_unit_0_register_file_0_r5[6]), .QN(), .CK(
      execution_unit_0_register_file_0_n_46), .D(
      execution_unit_0_register_file_0_n_53), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_139 (.ZN(
      execution_unit_0_register_file_0_n_105_133), .A1(
      execution_unit_0_register_file_0_n_45), .A2(
      execution_unit_0_register_file_0_r5[6]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_105_140 (.ZN(
      execution_unit_0_register_file_0_n_105_134), .A1(
      execution_unit_0_register_file_0_n_105_130), .A2(
      execution_unit_0_register_file_0_n_105_131), .A3(
      execution_unit_0_register_file_0_n_105_132), .A4(
      execution_unit_0_register_file_0_n_105_133));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_87_13 (.ZN(
      execution_unit_0_register_file_0_n_87_7), .A1(
      execution_unit_0_register_file_0_n_87_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[6]), .B1(
      execution_unit_0_register_file_0_r13_wr), .B2(execution_unit_0_alu_out[6]));
  INV_X1_LVT execution_unit_0_register_file_0_i_87_14 (.ZN(
      execution_unit_0_register_file_0_n_205), .A(
      execution_unit_0_register_file_0_n_87_7));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r13_reg[6] (.Q(
      execution_unit_0_register_file_0_r13[6]), .QN(), .CK(
      execution_unit_0_register_file_0_n_198), .D(
      execution_unit_0_register_file_0_n_205), .RN(
      execution_unit_0_register_file_0_n_8));
  AND2_X1_LVT execution_unit_0_register_file_0_i_105_141 (.ZN(
      execution_unit_0_register_file_0_n_105_135), .A1(
      execution_unit_0_register_file_0_n_197), .A2(
      execution_unit_0_register_file_0_r13[6]));
  NOR4_X1_LVT execution_unit_0_register_file_0_i_105_142 (.ZN(
      execution_unit_0_register_file_0_n_105_136), .A1(
      execution_unit_0_register_file_0_n_105_124), .A2(
      execution_unit_0_register_file_0_n_105_129), .A3(
      execution_unit_0_register_file_0_n_105_134), .A4(
      execution_unit_0_register_file_0_n_105_135));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_143 (.ZN(
      execution_unit_0_register_file_0_n_105_137), .A1(
      execution_unit_0_register_file_0_n_254), .A2(pc[6]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_101_13 (.ZN(
      execution_unit_0_register_file_0_n_101_7), .A1(
      execution_unit_0_register_file_0_n_101_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[6]), .B1(
      execution_unit_0_register_file_0_r15_wr), .B2(execution_unit_0_alu_out[6]));
  INV_X1_LVT execution_unit_0_register_file_0_i_101_14 (.ZN(
      execution_unit_0_register_file_0_n_243), .A(
      execution_unit_0_register_file_0_n_101_7));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r15_reg[6] (.Q(
      execution_unit_0_register_file_0_r15[6]), .QN(), .CK(
      execution_unit_0_register_file_0_n_236), .D(
      execution_unit_0_register_file_0_n_243), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_144 (.ZN(
      execution_unit_0_register_file_0_n_105_138), .A1(
      execution_unit_0_register_file_0_n_235), .A2(
      execution_unit_0_register_file_0_r15[6]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_94_13 (.ZN(
      execution_unit_0_register_file_0_n_94_7), .A1(
      execution_unit_0_register_file_0_n_94_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[6]), .B1(
      execution_unit_0_register_file_0_r14_wr), .B2(execution_unit_0_alu_out[6]));
  INV_X1_LVT execution_unit_0_register_file_0_i_94_14 (.ZN(
      execution_unit_0_register_file_0_n_224), .A(
      execution_unit_0_register_file_0_n_94_7));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r14_reg[6] (.Q(
      execution_unit_0_register_file_0_r14[6]), .QN(), .CK(
      execution_unit_0_register_file_0_n_217), .D(
      execution_unit_0_register_file_0_n_224), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_145 (.ZN(
      execution_unit_0_register_file_0_n_105_139), .A1(
      execution_unit_0_register_file_0_n_216), .A2(
      execution_unit_0_register_file_0_r14[6]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_105_146 (.ZN(
      execution_unit_0_reg_src[6]), .A1(
      execution_unit_0_register_file_0_n_105_136), .A2(
      execution_unit_0_register_file_0_n_105_137), .A3(
      execution_unit_0_register_file_0_n_105_138), .A4(
      execution_unit_0_register_file_0_n_105_139));
  HA_X1_LVT execution_unit_0_register_file_0_i_106_5 (.CO(
      execution_unit_0_register_file_0_n_106_4), .S(
      execution_unit_0_register_file_0_n_260), .A(execution_unit_0_reg_src[6]), 
      .B(execution_unit_0_register_file_0_n_106_3));
  HA_X1_LVT execution_unit_0_register_file_0_i_106_6 (.CO(
      execution_unit_0_register_file_0_n_106_5), .S(
      execution_unit_0_register_file_0_n_261), .A(execution_unit_0_reg_src[7]), 
      .B(execution_unit_0_register_file_0_n_106_4));
  AOI222_X1_LVT execution_unit_0_register_file_0_i_109_12 (.ZN(
      execution_unit_0_register_file_0_n_109_6), .A1(
      execution_unit_0_register_file_0_r1_wr), .A2(execution_unit_0_alu_out[7]), 
      .B1(execution_unit_0_register_file_0_n_272), .B2(eu_mab[7]), .C1(
      execution_unit_0_register_file_0_n_271), .C2(
      execution_unit_0_register_file_0_n_261));
  INV_X1_LVT execution_unit_0_register_file_0_i_109_13 (.ZN(
      execution_unit_0_register_file_0_n_279), .A(
      execution_unit_0_register_file_0_n_109_6));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r1_reg[7] (.Q(
      execution_unit_0_register_file_0_r1[7]), .QN(), .CK(
      execution_unit_0_register_file_0_n_270), .D(
      execution_unit_0_register_file_0_n_279), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_150 (.ZN(
      execution_unit_0_register_file_0_n_105_143), .A1(
      execution_unit_0_register_file_0_inst_src_in), .A2(
      execution_unit_0_register_file_0_r1[7]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_105_151 (.ZN(
      execution_unit_0_register_file_0_n_105_144), .A1(
      execution_unit_0_register_file_0_n_105_140), .A2(
      execution_unit_0_register_file_0_n_105_141), .A3(
      execution_unit_0_register_file_0_n_105_142), .A4(
      execution_unit_0_register_file_0_n_105_143));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_80_15 (.ZN(
      execution_unit_0_register_file_0_n_80_8), .A1(
      execution_unit_0_register_file_0_n_80_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[7]), .B1(
      execution_unit_0_register_file_0_r12_wr), .B2(execution_unit_0_alu_out[7]));
  INV_X1_LVT execution_unit_0_register_file_0_i_80_16 (.ZN(
      execution_unit_0_register_file_0_n_187), .A(
      execution_unit_0_register_file_0_n_80_8));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r12_reg[7] (.Q(
      execution_unit_0_register_file_0_r12[7]), .QN(), .CK(
      execution_unit_0_register_file_0_n_179), .D(
      execution_unit_0_register_file_0_n_187), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_152 (.ZN(
      execution_unit_0_register_file_0_n_105_145), .A1(
      execution_unit_0_register_file_0_n_178), .A2(
      execution_unit_0_register_file_0_r12[7]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_73_15 (.ZN(
      execution_unit_0_register_file_0_n_73_8), .A1(
      execution_unit_0_register_file_0_n_73_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[7]), .B1(
      execution_unit_0_register_file_0_r11_wr), .B2(execution_unit_0_alu_out[7]));
  INV_X1_LVT execution_unit_0_register_file_0_i_73_16 (.ZN(
      execution_unit_0_register_file_0_n_168), .A(
      execution_unit_0_register_file_0_n_73_8));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r11_reg[7] (.Q(
      execution_unit_0_register_file_0_r11[7]), .QN(), .CK(
      execution_unit_0_register_file_0_n_160), .D(
      execution_unit_0_register_file_0_n_168), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_153 (.ZN(
      execution_unit_0_register_file_0_n_105_146), .A1(
      execution_unit_0_register_file_0_n_159), .A2(
      execution_unit_0_register_file_0_r11[7]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_66_15 (.ZN(
      execution_unit_0_register_file_0_n_66_8), .A1(
      execution_unit_0_register_file_0_n_66_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[7]), .B1(
      execution_unit_0_register_file_0_r10_wr), .B2(execution_unit_0_alu_out[7]));
  INV_X1_LVT execution_unit_0_register_file_0_i_66_16 (.ZN(
      execution_unit_0_register_file_0_n_149), .A(
      execution_unit_0_register_file_0_n_66_8));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r10_reg[7] (.Q(
      execution_unit_0_register_file_0_r10[7]), .QN(), .CK(
      execution_unit_0_register_file_0_n_141), .D(
      execution_unit_0_register_file_0_n_149), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_154 (.ZN(
      execution_unit_0_register_file_0_n_105_147), .A1(
      execution_unit_0_register_file_0_n_140), .A2(
      execution_unit_0_register_file_0_r10[7]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_59_15 (.ZN(
      execution_unit_0_register_file_0_n_59_8), .A1(
      execution_unit_0_register_file_0_n_59_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[7]), .B1(
      execution_unit_0_register_file_0_r9_wr), .B2(execution_unit_0_alu_out[7]));
  INV_X1_LVT execution_unit_0_register_file_0_i_59_16 (.ZN(
      execution_unit_0_register_file_0_n_130), .A(
      execution_unit_0_register_file_0_n_59_8));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r9_reg[7] (.Q(
      execution_unit_0_register_file_0_r9[7]), .QN(), .CK(
      execution_unit_0_register_file_0_n_122), .D(
      execution_unit_0_register_file_0_n_130), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_155 (.ZN(
      execution_unit_0_register_file_0_n_105_148), .A1(
      execution_unit_0_register_file_0_n_121), .A2(
      execution_unit_0_register_file_0_r9[7]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_105_156 (.ZN(
      execution_unit_0_register_file_0_n_105_149), .A1(
      execution_unit_0_register_file_0_n_105_145), .A2(
      execution_unit_0_register_file_0_n_105_146), .A3(
      execution_unit_0_register_file_0_n_105_147), .A4(
      execution_unit_0_register_file_0_n_105_148));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_52_15 (.ZN(
      execution_unit_0_register_file_0_n_52_8), .A1(
      execution_unit_0_register_file_0_n_52_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[7]), .B1(
      execution_unit_0_register_file_0_r8_wr), .B2(execution_unit_0_alu_out[7]));
  INV_X1_LVT execution_unit_0_register_file_0_i_52_16 (.ZN(
      execution_unit_0_register_file_0_n_111), .A(
      execution_unit_0_register_file_0_n_52_8));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r8_reg[7] (.Q(
      execution_unit_0_register_file_0_r8[7]), .QN(), .CK(
      execution_unit_0_register_file_0_n_103), .D(
      execution_unit_0_register_file_0_n_111), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_157 (.ZN(
      execution_unit_0_register_file_0_n_105_150), .A1(
      execution_unit_0_register_file_0_n_102), .A2(
      execution_unit_0_register_file_0_r8[7]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_45_15 (.ZN(
      execution_unit_0_register_file_0_n_45_8), .A1(
      execution_unit_0_register_file_0_n_45_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[7]), .B1(
      execution_unit_0_register_file_0_r7_wr), .B2(execution_unit_0_alu_out[7]));
  INV_X1_LVT execution_unit_0_register_file_0_i_45_16 (.ZN(
      execution_unit_0_register_file_0_n_92), .A(
      execution_unit_0_register_file_0_n_45_8));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r7_reg[7] (.Q(
      execution_unit_0_register_file_0_r7[7]), .QN(), .CK(
      execution_unit_0_register_file_0_n_84), .D(
      execution_unit_0_register_file_0_n_92), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_158 (.ZN(
      execution_unit_0_register_file_0_n_105_151), .A1(
      execution_unit_0_register_file_0_n_83), .A2(
      execution_unit_0_register_file_0_r7[7]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_38_15 (.ZN(
      execution_unit_0_register_file_0_n_38_8), .A1(
      execution_unit_0_register_file_0_n_38_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[7]), .B1(
      execution_unit_0_register_file_0_r6_wr), .B2(execution_unit_0_alu_out[7]));
  INV_X1_LVT execution_unit_0_register_file_0_i_38_16 (.ZN(
      execution_unit_0_register_file_0_n_73), .A(
      execution_unit_0_register_file_0_n_38_8));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r6_reg[7] (.Q(
      execution_unit_0_register_file_0_r6[7]), .QN(), .CK(
      execution_unit_0_register_file_0_n_65), .D(
      execution_unit_0_register_file_0_n_73), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_159 (.ZN(
      execution_unit_0_register_file_0_n_105_152), .A1(
      execution_unit_0_register_file_0_n_64), .A2(
      execution_unit_0_register_file_0_r6[7]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_31_15 (.ZN(
      execution_unit_0_register_file_0_n_31_8), .A1(
      execution_unit_0_register_file_0_n_31_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[7]), .B1(
      execution_unit_0_register_file_0_r5_wr), .B2(execution_unit_0_alu_out[7]));
  INV_X1_LVT execution_unit_0_register_file_0_i_31_16 (.ZN(
      execution_unit_0_register_file_0_n_54), .A(
      execution_unit_0_register_file_0_n_31_8));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r5_reg[7] (.Q(
      execution_unit_0_register_file_0_r5[7]), .QN(), .CK(
      execution_unit_0_register_file_0_n_46), .D(
      execution_unit_0_register_file_0_n_54), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_160 (.ZN(
      execution_unit_0_register_file_0_n_105_153), .A1(
      execution_unit_0_register_file_0_n_45), .A2(
      execution_unit_0_register_file_0_r5[7]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_105_161 (.ZN(
      execution_unit_0_register_file_0_n_105_154), .A1(
      execution_unit_0_register_file_0_n_105_150), .A2(
      execution_unit_0_register_file_0_n_105_151), .A3(
      execution_unit_0_register_file_0_n_105_152), .A4(
      execution_unit_0_register_file_0_n_105_153));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_87_15 (.ZN(
      execution_unit_0_register_file_0_n_87_8), .A1(
      execution_unit_0_register_file_0_n_87_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[7]), .B1(
      execution_unit_0_register_file_0_r13_wr), .B2(execution_unit_0_alu_out[7]));
  INV_X1_LVT execution_unit_0_register_file_0_i_87_16 (.ZN(
      execution_unit_0_register_file_0_n_206), .A(
      execution_unit_0_register_file_0_n_87_8));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r13_reg[7] (.Q(
      execution_unit_0_register_file_0_r13[7]), .QN(), .CK(
      execution_unit_0_register_file_0_n_198), .D(
      execution_unit_0_register_file_0_n_206), .RN(
      execution_unit_0_register_file_0_n_8));
  AND2_X1_LVT execution_unit_0_register_file_0_i_105_162 (.ZN(
      execution_unit_0_register_file_0_n_105_155), .A1(
      execution_unit_0_register_file_0_n_197), .A2(
      execution_unit_0_register_file_0_r13[7]));
  NOR4_X1_LVT execution_unit_0_register_file_0_i_105_163 (.ZN(
      execution_unit_0_register_file_0_n_105_156), .A1(
      execution_unit_0_register_file_0_n_105_144), .A2(
      execution_unit_0_register_file_0_n_105_149), .A3(
      execution_unit_0_register_file_0_n_105_154), .A4(
      execution_unit_0_register_file_0_n_105_155));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_164 (.ZN(
      execution_unit_0_register_file_0_n_105_157), .A1(
      execution_unit_0_register_file_0_n_254), .A2(pc[7]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_101_15 (.ZN(
      execution_unit_0_register_file_0_n_101_8), .A1(
      execution_unit_0_register_file_0_n_101_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[7]), .B1(
      execution_unit_0_register_file_0_r15_wr), .B2(execution_unit_0_alu_out[7]));
  INV_X1_LVT execution_unit_0_register_file_0_i_101_16 (.ZN(
      execution_unit_0_register_file_0_n_244), .A(
      execution_unit_0_register_file_0_n_101_8));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r15_reg[7] (.Q(
      execution_unit_0_register_file_0_r15[7]), .QN(), .CK(
      execution_unit_0_register_file_0_n_236), .D(
      execution_unit_0_register_file_0_n_244), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_165 (.ZN(
      execution_unit_0_register_file_0_n_105_158), .A1(
      execution_unit_0_register_file_0_n_235), .A2(
      execution_unit_0_register_file_0_r15[7]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_94_15 (.ZN(
      execution_unit_0_register_file_0_n_94_8), .A1(
      execution_unit_0_register_file_0_n_94_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[7]), .B1(
      execution_unit_0_register_file_0_r14_wr), .B2(execution_unit_0_alu_out[7]));
  INV_X1_LVT execution_unit_0_register_file_0_i_94_16 (.ZN(
      execution_unit_0_register_file_0_n_225), .A(
      execution_unit_0_register_file_0_n_94_8));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r14_reg[7] (.Q(
      execution_unit_0_register_file_0_r14[7]), .QN(), .CK(
      execution_unit_0_register_file_0_n_217), .D(
      execution_unit_0_register_file_0_n_225), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_166 (.ZN(
      execution_unit_0_register_file_0_n_105_159), .A1(
      execution_unit_0_register_file_0_n_216), .A2(
      execution_unit_0_register_file_0_r14[7]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_105_167 (.ZN(
      execution_unit_0_reg_src[7]), .A1(
      execution_unit_0_register_file_0_n_105_156), .A2(
      execution_unit_0_register_file_0_n_105_157), .A3(
      execution_unit_0_register_file_0_n_105_158), .A4(
      execution_unit_0_register_file_0_n_105_159));
  HA_X1_LVT execution_unit_0_register_file_0_i_22_7 (.CO(
      execution_unit_0_register_file_0_n_22_7), .S(
      execution_unit_0_register_file_0_reg_incr_val[7]), .A(
      execution_unit_0_reg_src[7]), .B(execution_unit_0_register_file_0_n_22_6));
  HA_X1_LVT execution_unit_0_register_file_0_i_22_8 (.CO(
      execution_unit_0_register_file_0_n_22_8), .S(
      execution_unit_0_register_file_0_reg_incr_val[8]), .A(
      execution_unit_0_reg_src[8]), .B(execution_unit_0_register_file_0_n_22_7));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_24_17 (.ZN(
      execution_unit_0_register_file_0_n_24_9), .A1(
      execution_unit_0_register_file_0_n_24_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[8]), .B1(
      execution_unit_0_register_file_0_r4_wr), .B2(pc_sw[8]));
  INV_X1_LVT execution_unit_0_register_file_0_i_24_18 (.ZN(
      execution_unit_0_register_file_0_n_36), .A(
      execution_unit_0_register_file_0_n_24_9));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r4_reg[8] (.Q(
      execution_unit_0_register_file_0_r4[8]), .QN(), .CK(
      execution_unit_0_register_file_0_n_27), .D(
      execution_unit_0_register_file_0_n_36), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_168 (.ZN(
      execution_unit_0_register_file_0_n_105_160), .A1(
      execution_unit_0_register_file_0_n_24), .A2(
      execution_unit_0_register_file_0_r4[8]));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r3_reg[8] (.Q(
      execution_unit_0_register_file_0_r3[8]), .QN(), .CK(
      execution_unit_0_register_file_0_n_23), .D(pc_sw[8]), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_169 (.ZN(
      execution_unit_0_register_file_0_n_105_161), .A1(
      execution_unit_0_register_file_0_n_22), .A2(
      execution_unit_0_register_file_0_r3[8]));
  INV_X1_LVT execution_unit_0_register_file_0_i_5_16 (.ZN(
      execution_unit_0_register_file_0_n_5_13), .A(
      execution_unit_0_alu_stat_wr[3]));
  NAND3_X1_LVT execution_unit_0_register_file_0_i_5_17 (.ZN(
      execution_unit_0_register_file_0_n_5_14), .A1(
      execution_unit_0_register_file_0_n_5_0), .A2(
      execution_unit_0_register_file_0_n_5_13), .A3(execution_unit_0_status[3]));
  NAND3_X1_LVT execution_unit_0_register_file_0_i_5_18 (.ZN(
      execution_unit_0_register_file_0_n_5_15), .A1(
      execution_unit_0_register_file_0_n_5_13), .A2(
      execution_unit_0_register_file_0_r2_wr), .A3(pc_sw[8]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_5_19 (.ZN(
      execution_unit_0_register_file_0_n_5_16), .A1(execution_unit_0_alu_stat[3]), 
      .A2(execution_unit_0_alu_stat_wr[3]));
  NAND3_X1_LVT execution_unit_0_register_file_0_i_5_20 (.ZN(
      execution_unit_0_register_file_0_n_12), .A1(
      execution_unit_0_register_file_0_n_5_14), .A2(
      execution_unit_0_register_file_0_n_5_15), .A3(
      execution_unit_0_register_file_0_n_5_16));
  AND2_X1_LVT execution_unit_0_register_file_0_i_6_8 (.ZN(
      execution_unit_0_register_file_0_n_20), .A1(
      execution_unit_0_register_file_0_n_6_0), .A2(
      execution_unit_0_register_file_0_n_12));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r2_reg[8] (.Q(
      execution_unit_0_status[3]), .QN(), .CK(cpu_mclk), .D(
      execution_unit_0_register_file_0_n_20), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_170 (.ZN(
      execution_unit_0_register_file_0_n_105_162), .A1(
      execution_unit_0_register_file_0_n_21), .A2(execution_unit_0_status[3]));
  AOI222_X1_LVT execution_unit_0_register_file_0_i_109_14 (.ZN(
      execution_unit_0_register_file_0_n_109_7), .A1(
      execution_unit_0_register_file_0_r1_wr), .A2(pc_sw[8]), .B1(
      execution_unit_0_register_file_0_n_272), .B2(eu_mab[8]), .C1(
      execution_unit_0_register_file_0_n_271), .C2(
      execution_unit_0_register_file_0_n_262));
  INV_X1_LVT execution_unit_0_register_file_0_i_109_15 (.ZN(
      execution_unit_0_register_file_0_n_280), .A(
      execution_unit_0_register_file_0_n_109_7));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r1_reg[8] (.Q(
      execution_unit_0_register_file_0_r1[8]), .QN(), .CK(
      execution_unit_0_register_file_0_n_270), .D(
      execution_unit_0_register_file_0_n_280), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_171 (.ZN(
      execution_unit_0_register_file_0_n_105_163), .A1(
      execution_unit_0_register_file_0_inst_src_in), .A2(
      execution_unit_0_register_file_0_r1[8]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_105_172 (.ZN(
      execution_unit_0_register_file_0_n_105_164), .A1(
      execution_unit_0_register_file_0_n_105_160), .A2(
      execution_unit_0_register_file_0_n_105_161), .A3(
      execution_unit_0_register_file_0_n_105_162), .A4(
      execution_unit_0_register_file_0_n_105_163));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_80_17 (.ZN(
      execution_unit_0_register_file_0_n_80_9), .A1(
      execution_unit_0_register_file_0_n_80_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[8]), .B1(
      execution_unit_0_register_file_0_r12_wr), .B2(pc_sw[8]));
  INV_X1_LVT execution_unit_0_register_file_0_i_80_18 (.ZN(
      execution_unit_0_register_file_0_n_188), .A(
      execution_unit_0_register_file_0_n_80_9));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r12_reg[8] (.Q(
      execution_unit_0_register_file_0_r12[8]), .QN(), .CK(
      execution_unit_0_register_file_0_n_179), .D(
      execution_unit_0_register_file_0_n_188), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_173 (.ZN(
      execution_unit_0_register_file_0_n_105_165), .A1(
      execution_unit_0_register_file_0_n_178), .A2(
      execution_unit_0_register_file_0_r12[8]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_73_17 (.ZN(
      execution_unit_0_register_file_0_n_73_9), .A1(
      execution_unit_0_register_file_0_n_73_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[8]), .B1(
      execution_unit_0_register_file_0_r11_wr), .B2(pc_sw[8]));
  INV_X1_LVT execution_unit_0_register_file_0_i_73_18 (.ZN(
      execution_unit_0_register_file_0_n_169), .A(
      execution_unit_0_register_file_0_n_73_9));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r11_reg[8] (.Q(
      execution_unit_0_register_file_0_r11[8]), .QN(), .CK(
      execution_unit_0_register_file_0_n_160), .D(
      execution_unit_0_register_file_0_n_169), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_174 (.ZN(
      execution_unit_0_register_file_0_n_105_166), .A1(
      execution_unit_0_register_file_0_n_159), .A2(
      execution_unit_0_register_file_0_r11[8]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_66_17 (.ZN(
      execution_unit_0_register_file_0_n_66_9), .A1(
      execution_unit_0_register_file_0_n_66_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[8]), .B1(
      execution_unit_0_register_file_0_r10_wr), .B2(pc_sw[8]));
  INV_X1_LVT execution_unit_0_register_file_0_i_66_18 (.ZN(
      execution_unit_0_register_file_0_n_150), .A(
      execution_unit_0_register_file_0_n_66_9));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r10_reg[8] (.Q(
      execution_unit_0_register_file_0_r10[8]), .QN(), .CK(
      execution_unit_0_register_file_0_n_141), .D(
      execution_unit_0_register_file_0_n_150), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_175 (.ZN(
      execution_unit_0_register_file_0_n_105_167), .A1(
      execution_unit_0_register_file_0_n_140), .A2(
      execution_unit_0_register_file_0_r10[8]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_59_17 (.ZN(
      execution_unit_0_register_file_0_n_59_9), .A1(
      execution_unit_0_register_file_0_n_59_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[8]), .B1(
      execution_unit_0_register_file_0_r9_wr), .B2(pc_sw[8]));
  INV_X1_LVT execution_unit_0_register_file_0_i_59_18 (.ZN(
      execution_unit_0_register_file_0_n_131), .A(
      execution_unit_0_register_file_0_n_59_9));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r9_reg[8] (.Q(
      execution_unit_0_register_file_0_r9[8]), .QN(), .CK(
      execution_unit_0_register_file_0_n_122), .D(
      execution_unit_0_register_file_0_n_131), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_176 (.ZN(
      execution_unit_0_register_file_0_n_105_168), .A1(
      execution_unit_0_register_file_0_n_121), .A2(
      execution_unit_0_register_file_0_r9[8]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_105_177 (.ZN(
      execution_unit_0_register_file_0_n_105_169), .A1(
      execution_unit_0_register_file_0_n_105_165), .A2(
      execution_unit_0_register_file_0_n_105_166), .A3(
      execution_unit_0_register_file_0_n_105_167), .A4(
      execution_unit_0_register_file_0_n_105_168));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_52_17 (.ZN(
      execution_unit_0_register_file_0_n_52_9), .A1(
      execution_unit_0_register_file_0_n_52_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[8]), .B1(
      execution_unit_0_register_file_0_r8_wr), .B2(pc_sw[8]));
  INV_X1_LVT execution_unit_0_register_file_0_i_52_18 (.ZN(
      execution_unit_0_register_file_0_n_112), .A(
      execution_unit_0_register_file_0_n_52_9));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r8_reg[8] (.Q(
      execution_unit_0_register_file_0_r8[8]), .QN(), .CK(
      execution_unit_0_register_file_0_n_103), .D(
      execution_unit_0_register_file_0_n_112), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_178 (.ZN(
      execution_unit_0_register_file_0_n_105_170), .A1(
      execution_unit_0_register_file_0_n_102), .A2(
      execution_unit_0_register_file_0_r8[8]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_45_17 (.ZN(
      execution_unit_0_register_file_0_n_45_9), .A1(
      execution_unit_0_register_file_0_n_45_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[8]), .B1(
      execution_unit_0_register_file_0_r7_wr), .B2(pc_sw[8]));
  INV_X1_LVT execution_unit_0_register_file_0_i_45_18 (.ZN(
      execution_unit_0_register_file_0_n_93), .A(
      execution_unit_0_register_file_0_n_45_9));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r7_reg[8] (.Q(
      execution_unit_0_register_file_0_r7[8]), .QN(), .CK(
      execution_unit_0_register_file_0_n_84), .D(
      execution_unit_0_register_file_0_n_93), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_179 (.ZN(
      execution_unit_0_register_file_0_n_105_171), .A1(
      execution_unit_0_register_file_0_n_83), .A2(
      execution_unit_0_register_file_0_r7[8]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_38_17 (.ZN(
      execution_unit_0_register_file_0_n_38_9), .A1(
      execution_unit_0_register_file_0_n_38_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[8]), .B1(
      execution_unit_0_register_file_0_r6_wr), .B2(pc_sw[8]));
  INV_X1_LVT execution_unit_0_register_file_0_i_38_18 (.ZN(
      execution_unit_0_register_file_0_n_74), .A(
      execution_unit_0_register_file_0_n_38_9));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r6_reg[8] (.Q(
      execution_unit_0_register_file_0_r6[8]), .QN(), .CK(
      execution_unit_0_register_file_0_n_65), .D(
      execution_unit_0_register_file_0_n_74), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_180 (.ZN(
      execution_unit_0_register_file_0_n_105_172), .A1(
      execution_unit_0_register_file_0_n_64), .A2(
      execution_unit_0_register_file_0_r6[8]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_31_17 (.ZN(
      execution_unit_0_register_file_0_n_31_9), .A1(
      execution_unit_0_register_file_0_n_31_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[8]), .B1(
      execution_unit_0_register_file_0_r5_wr), .B2(pc_sw[8]));
  INV_X1_LVT execution_unit_0_register_file_0_i_31_18 (.ZN(
      execution_unit_0_register_file_0_n_55), .A(
      execution_unit_0_register_file_0_n_31_9));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r5_reg[8] (.Q(
      execution_unit_0_register_file_0_r5[8]), .QN(), .CK(
      execution_unit_0_register_file_0_n_46), .D(
      execution_unit_0_register_file_0_n_55), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_181 (.ZN(
      execution_unit_0_register_file_0_n_105_173), .A1(
      execution_unit_0_register_file_0_n_45), .A2(
      execution_unit_0_register_file_0_r5[8]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_105_182 (.ZN(
      execution_unit_0_register_file_0_n_105_174), .A1(
      execution_unit_0_register_file_0_n_105_170), .A2(
      execution_unit_0_register_file_0_n_105_171), .A3(
      execution_unit_0_register_file_0_n_105_172), .A4(
      execution_unit_0_register_file_0_n_105_173));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_87_17 (.ZN(
      execution_unit_0_register_file_0_n_87_9), .A1(
      execution_unit_0_register_file_0_n_87_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[8]), .B1(
      execution_unit_0_register_file_0_r13_wr), .B2(pc_sw[8]));
  INV_X1_LVT execution_unit_0_register_file_0_i_87_18 (.ZN(
      execution_unit_0_register_file_0_n_207), .A(
      execution_unit_0_register_file_0_n_87_9));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r13_reg[8] (.Q(
      execution_unit_0_register_file_0_r13[8]), .QN(), .CK(
      execution_unit_0_register_file_0_n_198), .D(
      execution_unit_0_register_file_0_n_207), .RN(
      execution_unit_0_register_file_0_n_8));
  AND2_X1_LVT execution_unit_0_register_file_0_i_105_183 (.ZN(
      execution_unit_0_register_file_0_n_105_175), .A1(
      execution_unit_0_register_file_0_n_197), .A2(
      execution_unit_0_register_file_0_r13[8]));
  NOR4_X1_LVT execution_unit_0_register_file_0_i_105_184 (.ZN(
      execution_unit_0_register_file_0_n_105_176), .A1(
      execution_unit_0_register_file_0_n_105_164), .A2(
      execution_unit_0_register_file_0_n_105_169), .A3(
      execution_unit_0_register_file_0_n_105_174), .A4(
      execution_unit_0_register_file_0_n_105_175));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_185 (.ZN(
      execution_unit_0_register_file_0_n_105_177), .A1(
      execution_unit_0_register_file_0_n_254), .A2(pc[8]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_101_17 (.ZN(
      execution_unit_0_register_file_0_n_101_9), .A1(
      execution_unit_0_register_file_0_n_101_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[8]), .B1(
      execution_unit_0_register_file_0_r15_wr), .B2(pc_sw[8]));
  INV_X1_LVT execution_unit_0_register_file_0_i_101_18 (.ZN(
      execution_unit_0_register_file_0_n_245), .A(
      execution_unit_0_register_file_0_n_101_9));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r15_reg[8] (.Q(
      execution_unit_0_register_file_0_r15[8]), .QN(), .CK(
      execution_unit_0_register_file_0_n_236), .D(
      execution_unit_0_register_file_0_n_245), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_186 (.ZN(
      execution_unit_0_register_file_0_n_105_178), .A1(
      execution_unit_0_register_file_0_n_235), .A2(
      execution_unit_0_register_file_0_r15[8]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_94_17 (.ZN(
      execution_unit_0_register_file_0_n_94_9), .A1(
      execution_unit_0_register_file_0_n_94_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[8]), .B1(
      execution_unit_0_register_file_0_r14_wr), .B2(pc_sw[8]));
  INV_X1_LVT execution_unit_0_register_file_0_i_94_18 (.ZN(
      execution_unit_0_register_file_0_n_226), .A(
      execution_unit_0_register_file_0_n_94_9));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r14_reg[8] (.Q(
      execution_unit_0_register_file_0_r14[8]), .QN(), .CK(
      execution_unit_0_register_file_0_n_217), .D(
      execution_unit_0_register_file_0_n_226), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_187 (.ZN(
      execution_unit_0_register_file_0_n_105_179), .A1(
      execution_unit_0_register_file_0_n_216), .A2(
      execution_unit_0_register_file_0_r14[8]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_105_188 (.ZN(
      execution_unit_0_reg_src[8]), .A1(
      execution_unit_0_register_file_0_n_105_176), .A2(
      execution_unit_0_register_file_0_n_105_177), .A3(
      execution_unit_0_register_file_0_n_105_178), .A4(
      execution_unit_0_register_file_0_n_105_179));
  HA_X1_LVT execution_unit_0_register_file_0_i_106_7 (.CO(
      execution_unit_0_register_file_0_n_106_6), .S(
      execution_unit_0_register_file_0_n_262), .A(execution_unit_0_reg_src[8]), 
      .B(execution_unit_0_register_file_0_n_106_5));
  HA_X1_LVT execution_unit_0_register_file_0_i_106_8 (.CO(
      execution_unit_0_register_file_0_n_106_7), .S(
      execution_unit_0_register_file_0_n_263), .A(execution_unit_0_reg_src[9]), 
      .B(execution_unit_0_register_file_0_n_106_6));
  AOI222_X1_LVT execution_unit_0_register_file_0_i_109_16 (.ZN(
      execution_unit_0_register_file_0_n_109_8), .A1(
      execution_unit_0_register_file_0_r1_wr), .A2(pc_sw[9]), .B1(
      execution_unit_0_register_file_0_n_272), .B2(eu_mab[9]), .C1(
      execution_unit_0_register_file_0_n_271), .C2(
      execution_unit_0_register_file_0_n_263));
  INV_X1_LVT execution_unit_0_register_file_0_i_109_17 (.ZN(
      execution_unit_0_register_file_0_n_281), .A(
      execution_unit_0_register_file_0_n_109_8));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r1_reg[9] (.Q(
      execution_unit_0_register_file_0_r1[9]), .QN(), .CK(
      execution_unit_0_register_file_0_n_270), .D(
      execution_unit_0_register_file_0_n_281), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_192 (.ZN(
      execution_unit_0_register_file_0_n_105_183), .A1(
      execution_unit_0_register_file_0_inst_src_in), .A2(
      execution_unit_0_register_file_0_r1[9]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_105_193 (.ZN(
      execution_unit_0_register_file_0_n_105_184), .A1(
      execution_unit_0_register_file_0_n_105_180), .A2(
      execution_unit_0_register_file_0_n_105_181), .A3(
      execution_unit_0_register_file_0_n_105_182), .A4(
      execution_unit_0_register_file_0_n_105_183));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_80_19 (.ZN(
      execution_unit_0_register_file_0_n_80_10), .A1(
      execution_unit_0_register_file_0_n_80_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[9]), .B1(
      execution_unit_0_register_file_0_r12_wr), .B2(pc_sw[9]));
  INV_X1_LVT execution_unit_0_register_file_0_i_80_20 (.ZN(
      execution_unit_0_register_file_0_n_189), .A(
      execution_unit_0_register_file_0_n_80_10));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r12_reg[9] (.Q(
      execution_unit_0_register_file_0_r12[9]), .QN(), .CK(
      execution_unit_0_register_file_0_n_179), .D(
      execution_unit_0_register_file_0_n_189), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_194 (.ZN(
      execution_unit_0_register_file_0_n_105_185), .A1(
      execution_unit_0_register_file_0_n_178), .A2(
      execution_unit_0_register_file_0_r12[9]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_73_19 (.ZN(
      execution_unit_0_register_file_0_n_73_10), .A1(
      execution_unit_0_register_file_0_n_73_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[9]), .B1(
      execution_unit_0_register_file_0_r11_wr), .B2(pc_sw[9]));
  INV_X1_LVT execution_unit_0_register_file_0_i_73_20 (.ZN(
      execution_unit_0_register_file_0_n_170), .A(
      execution_unit_0_register_file_0_n_73_10));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r11_reg[9] (.Q(
      execution_unit_0_register_file_0_r11[9]), .QN(), .CK(
      execution_unit_0_register_file_0_n_160), .D(
      execution_unit_0_register_file_0_n_170), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_195 (.ZN(
      execution_unit_0_register_file_0_n_105_186), .A1(
      execution_unit_0_register_file_0_n_159), .A2(
      execution_unit_0_register_file_0_r11[9]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_66_19 (.ZN(
      execution_unit_0_register_file_0_n_66_10), .A1(
      execution_unit_0_register_file_0_n_66_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[9]), .B1(
      execution_unit_0_register_file_0_r10_wr), .B2(pc_sw[9]));
  INV_X1_LVT execution_unit_0_register_file_0_i_66_20 (.ZN(
      execution_unit_0_register_file_0_n_151), .A(
      execution_unit_0_register_file_0_n_66_10));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r10_reg[9] (.Q(
      execution_unit_0_register_file_0_r10[9]), .QN(), .CK(
      execution_unit_0_register_file_0_n_141), .D(
      execution_unit_0_register_file_0_n_151), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_196 (.ZN(
      execution_unit_0_register_file_0_n_105_187), .A1(
      execution_unit_0_register_file_0_n_140), .A2(
      execution_unit_0_register_file_0_r10[9]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_59_19 (.ZN(
      execution_unit_0_register_file_0_n_59_10), .A1(
      execution_unit_0_register_file_0_n_59_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[9]), .B1(
      execution_unit_0_register_file_0_r9_wr), .B2(pc_sw[9]));
  INV_X1_LVT execution_unit_0_register_file_0_i_59_20 (.ZN(
      execution_unit_0_register_file_0_n_132), .A(
      execution_unit_0_register_file_0_n_59_10));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r9_reg[9] (.Q(
      execution_unit_0_register_file_0_r9[9]), .QN(), .CK(
      execution_unit_0_register_file_0_n_122), .D(
      execution_unit_0_register_file_0_n_132), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_197 (.ZN(
      execution_unit_0_register_file_0_n_105_188), .A1(
      execution_unit_0_register_file_0_n_121), .A2(
      execution_unit_0_register_file_0_r9[9]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_105_198 (.ZN(
      execution_unit_0_register_file_0_n_105_189), .A1(
      execution_unit_0_register_file_0_n_105_185), .A2(
      execution_unit_0_register_file_0_n_105_186), .A3(
      execution_unit_0_register_file_0_n_105_187), .A4(
      execution_unit_0_register_file_0_n_105_188));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_52_19 (.ZN(
      execution_unit_0_register_file_0_n_52_10), .A1(
      execution_unit_0_register_file_0_n_52_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[9]), .B1(
      execution_unit_0_register_file_0_r8_wr), .B2(pc_sw[9]));
  INV_X1_LVT execution_unit_0_register_file_0_i_52_20 (.ZN(
      execution_unit_0_register_file_0_n_113), .A(
      execution_unit_0_register_file_0_n_52_10));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r8_reg[9] (.Q(
      execution_unit_0_register_file_0_r8[9]), .QN(), .CK(
      execution_unit_0_register_file_0_n_103), .D(
      execution_unit_0_register_file_0_n_113), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_199 (.ZN(
      execution_unit_0_register_file_0_n_105_190), .A1(
      execution_unit_0_register_file_0_n_102), .A2(
      execution_unit_0_register_file_0_r8[9]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_45_19 (.ZN(
      execution_unit_0_register_file_0_n_45_10), .A1(
      execution_unit_0_register_file_0_n_45_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[9]), .B1(
      execution_unit_0_register_file_0_r7_wr), .B2(pc_sw[9]));
  INV_X1_LVT execution_unit_0_register_file_0_i_45_20 (.ZN(
      execution_unit_0_register_file_0_n_94), .A(
      execution_unit_0_register_file_0_n_45_10));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r7_reg[9] (.Q(
      execution_unit_0_register_file_0_r7[9]), .QN(), .CK(
      execution_unit_0_register_file_0_n_84), .D(
      execution_unit_0_register_file_0_n_94), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_200 (.ZN(
      execution_unit_0_register_file_0_n_105_191), .A1(
      execution_unit_0_register_file_0_n_83), .A2(
      execution_unit_0_register_file_0_r7[9]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_38_19 (.ZN(
      execution_unit_0_register_file_0_n_38_10), .A1(
      execution_unit_0_register_file_0_n_38_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[9]), .B1(
      execution_unit_0_register_file_0_r6_wr), .B2(pc_sw[9]));
  INV_X1_LVT execution_unit_0_register_file_0_i_38_20 (.ZN(
      execution_unit_0_register_file_0_n_75), .A(
      execution_unit_0_register_file_0_n_38_10));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r6_reg[9] (.Q(
      execution_unit_0_register_file_0_r6[9]), .QN(), .CK(
      execution_unit_0_register_file_0_n_65), .D(
      execution_unit_0_register_file_0_n_75), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_201 (.ZN(
      execution_unit_0_register_file_0_n_105_192), .A1(
      execution_unit_0_register_file_0_n_64), .A2(
      execution_unit_0_register_file_0_r6[9]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_31_19 (.ZN(
      execution_unit_0_register_file_0_n_31_10), .A1(
      execution_unit_0_register_file_0_n_31_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[9]), .B1(
      execution_unit_0_register_file_0_r5_wr), .B2(pc_sw[9]));
  INV_X1_LVT execution_unit_0_register_file_0_i_31_20 (.ZN(
      execution_unit_0_register_file_0_n_56), .A(
      execution_unit_0_register_file_0_n_31_10));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r5_reg[9] (.Q(
      execution_unit_0_register_file_0_r5[9]), .QN(), .CK(
      execution_unit_0_register_file_0_n_46), .D(
      execution_unit_0_register_file_0_n_56), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_202 (.ZN(
      execution_unit_0_register_file_0_n_105_193), .A1(
      execution_unit_0_register_file_0_n_45), .A2(
      execution_unit_0_register_file_0_r5[9]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_105_203 (.ZN(
      execution_unit_0_register_file_0_n_105_194), .A1(
      execution_unit_0_register_file_0_n_105_190), .A2(
      execution_unit_0_register_file_0_n_105_191), .A3(
      execution_unit_0_register_file_0_n_105_192), .A4(
      execution_unit_0_register_file_0_n_105_193));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_87_19 (.ZN(
      execution_unit_0_register_file_0_n_87_10), .A1(
      execution_unit_0_register_file_0_n_87_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[9]), .B1(
      execution_unit_0_register_file_0_r13_wr), .B2(pc_sw[9]));
  INV_X1_LVT execution_unit_0_register_file_0_i_87_20 (.ZN(
      execution_unit_0_register_file_0_n_208), .A(
      execution_unit_0_register_file_0_n_87_10));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r13_reg[9] (.Q(
      execution_unit_0_register_file_0_r13[9]), .QN(), .CK(
      execution_unit_0_register_file_0_n_198), .D(
      execution_unit_0_register_file_0_n_208), .RN(
      execution_unit_0_register_file_0_n_8));
  AND2_X1_LVT execution_unit_0_register_file_0_i_105_204 (.ZN(
      execution_unit_0_register_file_0_n_105_195), .A1(
      execution_unit_0_register_file_0_n_197), .A2(
      execution_unit_0_register_file_0_r13[9]));
  NOR4_X1_LVT execution_unit_0_register_file_0_i_105_205 (.ZN(
      execution_unit_0_register_file_0_n_105_196), .A1(
      execution_unit_0_register_file_0_n_105_184), .A2(
      execution_unit_0_register_file_0_n_105_189), .A3(
      execution_unit_0_register_file_0_n_105_194), .A4(
      execution_unit_0_register_file_0_n_105_195));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_206 (.ZN(
      execution_unit_0_register_file_0_n_105_197), .A1(
      execution_unit_0_register_file_0_n_254), .A2(pc[9]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_101_19 (.ZN(
      execution_unit_0_register_file_0_n_101_10), .A1(
      execution_unit_0_register_file_0_n_101_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[9]), .B1(
      execution_unit_0_register_file_0_r15_wr), .B2(pc_sw[9]));
  INV_X1_LVT execution_unit_0_register_file_0_i_101_20 (.ZN(
      execution_unit_0_register_file_0_n_246), .A(
      execution_unit_0_register_file_0_n_101_10));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r15_reg[9] (.Q(
      execution_unit_0_register_file_0_r15[9]), .QN(), .CK(
      execution_unit_0_register_file_0_n_236), .D(
      execution_unit_0_register_file_0_n_246), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_207 (.ZN(
      execution_unit_0_register_file_0_n_105_198), .A1(
      execution_unit_0_register_file_0_n_235), .A2(
      execution_unit_0_register_file_0_r15[9]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_94_19 (.ZN(
      execution_unit_0_register_file_0_n_94_10), .A1(
      execution_unit_0_register_file_0_n_94_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[9]), .B1(
      execution_unit_0_register_file_0_r14_wr), .B2(pc_sw[9]));
  INV_X1_LVT execution_unit_0_register_file_0_i_94_20 (.ZN(
      execution_unit_0_register_file_0_n_227), .A(
      execution_unit_0_register_file_0_n_94_10));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r14_reg[9] (.Q(
      execution_unit_0_register_file_0_r14[9]), .QN(), .CK(
      execution_unit_0_register_file_0_n_217), .D(
      execution_unit_0_register_file_0_n_227), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_208 (.ZN(
      execution_unit_0_register_file_0_n_105_199), .A1(
      execution_unit_0_register_file_0_n_216), .A2(
      execution_unit_0_register_file_0_r14[9]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_105_209 (.ZN(
      execution_unit_0_reg_src[9]), .A1(
      execution_unit_0_register_file_0_n_105_196), .A2(
      execution_unit_0_register_file_0_n_105_197), .A3(
      execution_unit_0_register_file_0_n_105_198), .A4(
      execution_unit_0_register_file_0_n_105_199));
  HA_X1_LVT execution_unit_0_register_file_0_i_22_9 (.CO(
      execution_unit_0_register_file_0_n_22_9), .S(
      execution_unit_0_register_file_0_reg_incr_val[9]), .A(
      execution_unit_0_reg_src[9]), .B(execution_unit_0_register_file_0_n_22_8));
  HA_X1_LVT execution_unit_0_register_file_0_i_22_10 (.CO(
      execution_unit_0_register_file_0_n_22_10), .S(
      execution_unit_0_register_file_0_reg_incr_val[10]), .A(
      execution_unit_0_reg_src[10]), .B(execution_unit_0_register_file_0_n_22_9));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_24_21 (.ZN(
      execution_unit_0_register_file_0_n_24_11), .A1(
      execution_unit_0_register_file_0_n_24_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[10]), .B1(
      execution_unit_0_register_file_0_r4_wr), .B2(pc_sw[10]));
  INV_X1_LVT execution_unit_0_register_file_0_i_24_22 (.ZN(
      execution_unit_0_register_file_0_n_38), .A(
      execution_unit_0_register_file_0_n_24_11));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r4_reg[10] (.Q(
      execution_unit_0_register_file_0_r4[10]), .QN(), .CK(
      execution_unit_0_register_file_0_n_27), .D(
      execution_unit_0_register_file_0_n_38), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_210 (.ZN(
      execution_unit_0_register_file_0_n_105_200), .A1(
      execution_unit_0_register_file_0_n_24), .A2(
      execution_unit_0_register_file_0_r4[10]));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r3_reg[10] (.Q(
      execution_unit_0_register_file_0_r3[10]), .QN(), .CK(
      execution_unit_0_register_file_0_n_23), .D(pc_sw[10]), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_211 (.ZN(
      execution_unit_0_register_file_0_n_105_201), .A1(
      execution_unit_0_register_file_0_n_22), .A2(
      execution_unit_0_register_file_0_r3[10]));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r2_reg[10] (.Q(
      execution_unit_0_register_file_0_n_5), .QN(), .CK(cpu_mclk), .D(1'b0), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_212 (.ZN(
      execution_unit_0_register_file_0_n_105_202), .A1(
      execution_unit_0_register_file_0_n_21), .A2(
      execution_unit_0_register_file_0_n_5));
  AOI222_X1_LVT execution_unit_0_register_file_0_i_109_18 (.ZN(
      execution_unit_0_register_file_0_n_109_9), .A1(
      execution_unit_0_register_file_0_r1_wr), .A2(pc_sw[10]), .B1(
      execution_unit_0_register_file_0_n_272), .B2(eu_mab[10]), .C1(
      execution_unit_0_register_file_0_n_271), .C2(
      execution_unit_0_register_file_0_n_264));
  INV_X1_LVT execution_unit_0_register_file_0_i_109_19 (.ZN(
      execution_unit_0_register_file_0_n_282), .A(
      execution_unit_0_register_file_0_n_109_9));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r1_reg[10] (.Q(
      execution_unit_0_register_file_0_r1[10]), .QN(), .CK(
      execution_unit_0_register_file_0_n_270), .D(
      execution_unit_0_register_file_0_n_282), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_213 (.ZN(
      execution_unit_0_register_file_0_n_105_203), .A1(
      execution_unit_0_register_file_0_inst_src_in), .A2(
      execution_unit_0_register_file_0_r1[10]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_105_214 (.ZN(
      execution_unit_0_register_file_0_n_105_204), .A1(
      execution_unit_0_register_file_0_n_105_200), .A2(
      execution_unit_0_register_file_0_n_105_201), .A3(
      execution_unit_0_register_file_0_n_105_202), .A4(
      execution_unit_0_register_file_0_n_105_203));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_80_21 (.ZN(
      execution_unit_0_register_file_0_n_80_11), .A1(
      execution_unit_0_register_file_0_n_80_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[10]), .B1(
      execution_unit_0_register_file_0_r12_wr), .B2(pc_sw[10]));
  INV_X1_LVT execution_unit_0_register_file_0_i_80_22 (.ZN(
      execution_unit_0_register_file_0_n_190), .A(
      execution_unit_0_register_file_0_n_80_11));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r12_reg[10] (.Q(
      execution_unit_0_register_file_0_r12[10]), .QN(), .CK(
      execution_unit_0_register_file_0_n_179), .D(
      execution_unit_0_register_file_0_n_190), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_215 (.ZN(
      execution_unit_0_register_file_0_n_105_205), .A1(
      execution_unit_0_register_file_0_n_178), .A2(
      execution_unit_0_register_file_0_r12[10]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_73_21 (.ZN(
      execution_unit_0_register_file_0_n_73_11), .A1(
      execution_unit_0_register_file_0_n_73_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[10]), .B1(
      execution_unit_0_register_file_0_r11_wr), .B2(pc_sw[10]));
  INV_X1_LVT execution_unit_0_register_file_0_i_73_22 (.ZN(
      execution_unit_0_register_file_0_n_171), .A(
      execution_unit_0_register_file_0_n_73_11));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r11_reg[10] (.Q(
      execution_unit_0_register_file_0_r11[10]), .QN(), .CK(
      execution_unit_0_register_file_0_n_160), .D(
      execution_unit_0_register_file_0_n_171), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_216 (.ZN(
      execution_unit_0_register_file_0_n_105_206), .A1(
      execution_unit_0_register_file_0_n_159), .A2(
      execution_unit_0_register_file_0_r11[10]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_66_21 (.ZN(
      execution_unit_0_register_file_0_n_66_11), .A1(
      execution_unit_0_register_file_0_n_66_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[10]), .B1(
      execution_unit_0_register_file_0_r10_wr), .B2(pc_sw[10]));
  INV_X1_LVT execution_unit_0_register_file_0_i_66_22 (.ZN(
      execution_unit_0_register_file_0_n_152), .A(
      execution_unit_0_register_file_0_n_66_11));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r10_reg[10] (.Q(
      execution_unit_0_register_file_0_r10[10]), .QN(), .CK(
      execution_unit_0_register_file_0_n_141), .D(
      execution_unit_0_register_file_0_n_152), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_217 (.ZN(
      execution_unit_0_register_file_0_n_105_207), .A1(
      execution_unit_0_register_file_0_n_140), .A2(
      execution_unit_0_register_file_0_r10[10]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_59_21 (.ZN(
      execution_unit_0_register_file_0_n_59_11), .A1(
      execution_unit_0_register_file_0_n_59_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[10]), .B1(
      execution_unit_0_register_file_0_r9_wr), .B2(pc_sw[10]));
  INV_X1_LVT execution_unit_0_register_file_0_i_59_22 (.ZN(
      execution_unit_0_register_file_0_n_133), .A(
      execution_unit_0_register_file_0_n_59_11));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r9_reg[10] (.Q(
      execution_unit_0_register_file_0_r9[10]), .QN(), .CK(
      execution_unit_0_register_file_0_n_122), .D(
      execution_unit_0_register_file_0_n_133), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_218 (.ZN(
      execution_unit_0_register_file_0_n_105_208), .A1(
      execution_unit_0_register_file_0_n_121), .A2(
      execution_unit_0_register_file_0_r9[10]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_105_219 (.ZN(
      execution_unit_0_register_file_0_n_105_209), .A1(
      execution_unit_0_register_file_0_n_105_205), .A2(
      execution_unit_0_register_file_0_n_105_206), .A3(
      execution_unit_0_register_file_0_n_105_207), .A4(
      execution_unit_0_register_file_0_n_105_208));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_52_21 (.ZN(
      execution_unit_0_register_file_0_n_52_11), .A1(
      execution_unit_0_register_file_0_n_52_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[10]), .B1(
      execution_unit_0_register_file_0_r8_wr), .B2(pc_sw[10]));
  INV_X1_LVT execution_unit_0_register_file_0_i_52_22 (.ZN(
      execution_unit_0_register_file_0_n_114), .A(
      execution_unit_0_register_file_0_n_52_11));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r8_reg[10] (.Q(
      execution_unit_0_register_file_0_r8[10]), .QN(), .CK(
      execution_unit_0_register_file_0_n_103), .D(
      execution_unit_0_register_file_0_n_114), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_220 (.ZN(
      execution_unit_0_register_file_0_n_105_210), .A1(
      execution_unit_0_register_file_0_n_102), .A2(
      execution_unit_0_register_file_0_r8[10]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_45_21 (.ZN(
      execution_unit_0_register_file_0_n_45_11), .A1(
      execution_unit_0_register_file_0_n_45_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[10]), .B1(
      execution_unit_0_register_file_0_r7_wr), .B2(pc_sw[10]));
  INV_X1_LVT execution_unit_0_register_file_0_i_45_22 (.ZN(
      execution_unit_0_register_file_0_n_95), .A(
      execution_unit_0_register_file_0_n_45_11));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r7_reg[10] (.Q(
      execution_unit_0_register_file_0_r7[10]), .QN(), .CK(
      execution_unit_0_register_file_0_n_84), .D(
      execution_unit_0_register_file_0_n_95), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_221 (.ZN(
      execution_unit_0_register_file_0_n_105_211), .A1(
      execution_unit_0_register_file_0_n_83), .A2(
      execution_unit_0_register_file_0_r7[10]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_38_21 (.ZN(
      execution_unit_0_register_file_0_n_38_11), .A1(
      execution_unit_0_register_file_0_n_38_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[10]), .B1(
      execution_unit_0_register_file_0_r6_wr), .B2(pc_sw[10]));
  INV_X1_LVT execution_unit_0_register_file_0_i_38_22 (.ZN(
      execution_unit_0_register_file_0_n_76), .A(
      execution_unit_0_register_file_0_n_38_11));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r6_reg[10] (.Q(
      execution_unit_0_register_file_0_r6[10]), .QN(), .CK(
      execution_unit_0_register_file_0_n_65), .D(
      execution_unit_0_register_file_0_n_76), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_222 (.ZN(
      execution_unit_0_register_file_0_n_105_212), .A1(
      execution_unit_0_register_file_0_n_64), .A2(
      execution_unit_0_register_file_0_r6[10]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_31_21 (.ZN(
      execution_unit_0_register_file_0_n_31_11), .A1(
      execution_unit_0_register_file_0_n_31_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[10]), .B1(
      execution_unit_0_register_file_0_r5_wr), .B2(pc_sw[10]));
  INV_X1_LVT execution_unit_0_register_file_0_i_31_22 (.ZN(
      execution_unit_0_register_file_0_n_57), .A(
      execution_unit_0_register_file_0_n_31_11));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r5_reg[10] (.Q(
      execution_unit_0_register_file_0_r5[10]), .QN(), .CK(
      execution_unit_0_register_file_0_n_46), .D(
      execution_unit_0_register_file_0_n_57), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_223 (.ZN(
      execution_unit_0_register_file_0_n_105_213), .A1(
      execution_unit_0_register_file_0_n_45), .A2(
      execution_unit_0_register_file_0_r5[10]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_105_224 (.ZN(
      execution_unit_0_register_file_0_n_105_214), .A1(
      execution_unit_0_register_file_0_n_105_210), .A2(
      execution_unit_0_register_file_0_n_105_211), .A3(
      execution_unit_0_register_file_0_n_105_212), .A4(
      execution_unit_0_register_file_0_n_105_213));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_87_21 (.ZN(
      execution_unit_0_register_file_0_n_87_11), .A1(
      execution_unit_0_register_file_0_n_87_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[10]), .B1(
      execution_unit_0_register_file_0_r13_wr), .B2(pc_sw[10]));
  INV_X1_LVT execution_unit_0_register_file_0_i_87_22 (.ZN(
      execution_unit_0_register_file_0_n_209), .A(
      execution_unit_0_register_file_0_n_87_11));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r13_reg[10] (.Q(
      execution_unit_0_register_file_0_r13[10]), .QN(), .CK(
      execution_unit_0_register_file_0_n_198), .D(
      execution_unit_0_register_file_0_n_209), .RN(
      execution_unit_0_register_file_0_n_8));
  AND2_X1_LVT execution_unit_0_register_file_0_i_105_225 (.ZN(
      execution_unit_0_register_file_0_n_105_215), .A1(
      execution_unit_0_register_file_0_n_197), .A2(
      execution_unit_0_register_file_0_r13[10]));
  NOR4_X1_LVT execution_unit_0_register_file_0_i_105_226 (.ZN(
      execution_unit_0_register_file_0_n_105_216), .A1(
      execution_unit_0_register_file_0_n_105_204), .A2(
      execution_unit_0_register_file_0_n_105_209), .A3(
      execution_unit_0_register_file_0_n_105_214), .A4(
      execution_unit_0_register_file_0_n_105_215));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_227 (.ZN(
      execution_unit_0_register_file_0_n_105_217), .A1(
      execution_unit_0_register_file_0_n_254), .A2(pc[10]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_101_21 (.ZN(
      execution_unit_0_register_file_0_n_101_11), .A1(
      execution_unit_0_register_file_0_n_101_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[10]), .B1(
      execution_unit_0_register_file_0_r15_wr), .B2(pc_sw[10]));
  INV_X1_LVT execution_unit_0_register_file_0_i_101_22 (.ZN(
      execution_unit_0_register_file_0_n_247), .A(
      execution_unit_0_register_file_0_n_101_11));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r15_reg[10] (.Q(
      execution_unit_0_register_file_0_r15[10]), .QN(), .CK(
      execution_unit_0_register_file_0_n_236), .D(
      execution_unit_0_register_file_0_n_247), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_228 (.ZN(
      execution_unit_0_register_file_0_n_105_218), .A1(
      execution_unit_0_register_file_0_n_235), .A2(
      execution_unit_0_register_file_0_r15[10]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_94_21 (.ZN(
      execution_unit_0_register_file_0_n_94_11), .A1(
      execution_unit_0_register_file_0_n_94_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[10]), .B1(
      execution_unit_0_register_file_0_r14_wr), .B2(pc_sw[10]));
  INV_X1_LVT execution_unit_0_register_file_0_i_94_22 (.ZN(
      execution_unit_0_register_file_0_n_228), .A(
      execution_unit_0_register_file_0_n_94_11));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r14_reg[10] (.Q(
      execution_unit_0_register_file_0_r14[10]), .QN(), .CK(
      execution_unit_0_register_file_0_n_217), .D(
      execution_unit_0_register_file_0_n_228), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_229 (.ZN(
      execution_unit_0_register_file_0_n_105_219), .A1(
      execution_unit_0_register_file_0_n_216), .A2(
      execution_unit_0_register_file_0_r14[10]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_105_230 (.ZN(
      execution_unit_0_reg_src[10]), .A1(
      execution_unit_0_register_file_0_n_105_216), .A2(
      execution_unit_0_register_file_0_n_105_217), .A3(
      execution_unit_0_register_file_0_n_105_218), .A4(
      execution_unit_0_register_file_0_n_105_219));
  HA_X1_LVT execution_unit_0_register_file_0_i_106_9 (.CO(
      execution_unit_0_register_file_0_n_106_8), .S(
      execution_unit_0_register_file_0_n_264), .A(execution_unit_0_reg_src[10]), 
      .B(execution_unit_0_register_file_0_n_106_7));
  HA_X1_LVT execution_unit_0_register_file_0_i_106_10 (.CO(
      execution_unit_0_register_file_0_n_106_9), .S(
      execution_unit_0_register_file_0_n_265), .A(execution_unit_0_reg_src[11]), 
      .B(execution_unit_0_register_file_0_n_106_8));
  AOI222_X1_LVT execution_unit_0_register_file_0_i_109_20 (.ZN(
      execution_unit_0_register_file_0_n_109_10), .A1(
      execution_unit_0_register_file_0_r1_wr), .A2(pc_sw[11]), .B1(
      execution_unit_0_register_file_0_n_272), .B2(eu_mab[11]), .C1(
      execution_unit_0_register_file_0_n_271), .C2(
      execution_unit_0_register_file_0_n_265));
  INV_X1_LVT execution_unit_0_register_file_0_i_109_21 (.ZN(
      execution_unit_0_register_file_0_n_283), .A(
      execution_unit_0_register_file_0_n_109_10));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r1_reg[11] (.Q(
      execution_unit_0_register_file_0_r1[11]), .QN(), .CK(
      execution_unit_0_register_file_0_n_270), .D(
      execution_unit_0_register_file_0_n_283), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_234 (.ZN(
      execution_unit_0_register_file_0_n_105_223), .A1(
      execution_unit_0_register_file_0_inst_src_in), .A2(
      execution_unit_0_register_file_0_r1[11]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_105_235 (.ZN(
      execution_unit_0_register_file_0_n_105_224), .A1(
      execution_unit_0_register_file_0_n_105_220), .A2(
      execution_unit_0_register_file_0_n_105_221), .A3(
      execution_unit_0_register_file_0_n_105_222), .A4(
      execution_unit_0_register_file_0_n_105_223));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_80_23 (.ZN(
      execution_unit_0_register_file_0_n_80_12), .A1(
      execution_unit_0_register_file_0_n_80_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[11]), .B1(
      execution_unit_0_register_file_0_r12_wr), .B2(pc_sw[11]));
  INV_X1_LVT execution_unit_0_register_file_0_i_80_24 (.ZN(
      execution_unit_0_register_file_0_n_191), .A(
      execution_unit_0_register_file_0_n_80_12));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r12_reg[11] (.Q(
      execution_unit_0_register_file_0_r12[11]), .QN(), .CK(
      execution_unit_0_register_file_0_n_179), .D(
      execution_unit_0_register_file_0_n_191), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_236 (.ZN(
      execution_unit_0_register_file_0_n_105_225), .A1(
      execution_unit_0_register_file_0_n_178), .A2(
      execution_unit_0_register_file_0_r12[11]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_73_23 (.ZN(
      execution_unit_0_register_file_0_n_73_12), .A1(
      execution_unit_0_register_file_0_n_73_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[11]), .B1(
      execution_unit_0_register_file_0_r11_wr), .B2(pc_sw[11]));
  INV_X1_LVT execution_unit_0_register_file_0_i_73_24 (.ZN(
      execution_unit_0_register_file_0_n_172), .A(
      execution_unit_0_register_file_0_n_73_12));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r11_reg[11] (.Q(
      execution_unit_0_register_file_0_r11[11]), .QN(), .CK(
      execution_unit_0_register_file_0_n_160), .D(
      execution_unit_0_register_file_0_n_172), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_237 (.ZN(
      execution_unit_0_register_file_0_n_105_226), .A1(
      execution_unit_0_register_file_0_n_159), .A2(
      execution_unit_0_register_file_0_r11[11]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_66_23 (.ZN(
      execution_unit_0_register_file_0_n_66_12), .A1(
      execution_unit_0_register_file_0_n_66_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[11]), .B1(
      execution_unit_0_register_file_0_r10_wr), .B2(pc_sw[11]));
  INV_X1_LVT execution_unit_0_register_file_0_i_66_24 (.ZN(
      execution_unit_0_register_file_0_n_153), .A(
      execution_unit_0_register_file_0_n_66_12));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r10_reg[11] (.Q(
      execution_unit_0_register_file_0_r10[11]), .QN(), .CK(
      execution_unit_0_register_file_0_n_141), .D(
      execution_unit_0_register_file_0_n_153), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_238 (.ZN(
      execution_unit_0_register_file_0_n_105_227), .A1(
      execution_unit_0_register_file_0_n_140), .A2(
      execution_unit_0_register_file_0_r10[11]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_59_23 (.ZN(
      execution_unit_0_register_file_0_n_59_12), .A1(
      execution_unit_0_register_file_0_n_59_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[11]), .B1(
      execution_unit_0_register_file_0_r9_wr), .B2(pc_sw[11]));
  INV_X1_LVT execution_unit_0_register_file_0_i_59_24 (.ZN(
      execution_unit_0_register_file_0_n_134), .A(
      execution_unit_0_register_file_0_n_59_12));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r9_reg[11] (.Q(
      execution_unit_0_register_file_0_r9[11]), .QN(), .CK(
      execution_unit_0_register_file_0_n_122), .D(
      execution_unit_0_register_file_0_n_134), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_239 (.ZN(
      execution_unit_0_register_file_0_n_105_228), .A1(
      execution_unit_0_register_file_0_n_121), .A2(
      execution_unit_0_register_file_0_r9[11]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_105_240 (.ZN(
      execution_unit_0_register_file_0_n_105_229), .A1(
      execution_unit_0_register_file_0_n_105_225), .A2(
      execution_unit_0_register_file_0_n_105_226), .A3(
      execution_unit_0_register_file_0_n_105_227), .A4(
      execution_unit_0_register_file_0_n_105_228));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_52_23 (.ZN(
      execution_unit_0_register_file_0_n_52_12), .A1(
      execution_unit_0_register_file_0_n_52_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[11]), .B1(
      execution_unit_0_register_file_0_r8_wr), .B2(pc_sw[11]));
  INV_X1_LVT execution_unit_0_register_file_0_i_52_24 (.ZN(
      execution_unit_0_register_file_0_n_115), .A(
      execution_unit_0_register_file_0_n_52_12));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r8_reg[11] (.Q(
      execution_unit_0_register_file_0_r8[11]), .QN(), .CK(
      execution_unit_0_register_file_0_n_103), .D(
      execution_unit_0_register_file_0_n_115), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_241 (.ZN(
      execution_unit_0_register_file_0_n_105_230), .A1(
      execution_unit_0_register_file_0_n_102), .A2(
      execution_unit_0_register_file_0_r8[11]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_45_23 (.ZN(
      execution_unit_0_register_file_0_n_45_12), .A1(
      execution_unit_0_register_file_0_n_45_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[11]), .B1(
      execution_unit_0_register_file_0_r7_wr), .B2(pc_sw[11]));
  INV_X1_LVT execution_unit_0_register_file_0_i_45_24 (.ZN(
      execution_unit_0_register_file_0_n_96), .A(
      execution_unit_0_register_file_0_n_45_12));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r7_reg[11] (.Q(
      execution_unit_0_register_file_0_r7[11]), .QN(), .CK(
      execution_unit_0_register_file_0_n_84), .D(
      execution_unit_0_register_file_0_n_96), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_242 (.ZN(
      execution_unit_0_register_file_0_n_105_231), .A1(
      execution_unit_0_register_file_0_n_83), .A2(
      execution_unit_0_register_file_0_r7[11]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_38_23 (.ZN(
      execution_unit_0_register_file_0_n_38_12), .A1(
      execution_unit_0_register_file_0_n_38_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[11]), .B1(
      execution_unit_0_register_file_0_r6_wr), .B2(pc_sw[11]));
  INV_X1_LVT execution_unit_0_register_file_0_i_38_24 (.ZN(
      execution_unit_0_register_file_0_n_77), .A(
      execution_unit_0_register_file_0_n_38_12));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r6_reg[11] (.Q(
      execution_unit_0_register_file_0_r6[11]), .QN(), .CK(
      execution_unit_0_register_file_0_n_65), .D(
      execution_unit_0_register_file_0_n_77), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_243 (.ZN(
      execution_unit_0_register_file_0_n_105_232), .A1(
      execution_unit_0_register_file_0_n_64), .A2(
      execution_unit_0_register_file_0_r6[11]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_31_23 (.ZN(
      execution_unit_0_register_file_0_n_31_12), .A1(
      execution_unit_0_register_file_0_n_31_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[11]), .B1(
      execution_unit_0_register_file_0_r5_wr), .B2(pc_sw[11]));
  INV_X1_LVT execution_unit_0_register_file_0_i_31_24 (.ZN(
      execution_unit_0_register_file_0_n_58), .A(
      execution_unit_0_register_file_0_n_31_12));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r5_reg[11] (.Q(
      execution_unit_0_register_file_0_r5[11]), .QN(), .CK(
      execution_unit_0_register_file_0_n_46), .D(
      execution_unit_0_register_file_0_n_58), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_244 (.ZN(
      execution_unit_0_register_file_0_n_105_233), .A1(
      execution_unit_0_register_file_0_n_45), .A2(
      execution_unit_0_register_file_0_r5[11]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_105_245 (.ZN(
      execution_unit_0_register_file_0_n_105_234), .A1(
      execution_unit_0_register_file_0_n_105_230), .A2(
      execution_unit_0_register_file_0_n_105_231), .A3(
      execution_unit_0_register_file_0_n_105_232), .A4(
      execution_unit_0_register_file_0_n_105_233));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_87_23 (.ZN(
      execution_unit_0_register_file_0_n_87_12), .A1(
      execution_unit_0_register_file_0_n_87_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[11]), .B1(
      execution_unit_0_register_file_0_r13_wr), .B2(pc_sw[11]));
  INV_X1_LVT execution_unit_0_register_file_0_i_87_24 (.ZN(
      execution_unit_0_register_file_0_n_210), .A(
      execution_unit_0_register_file_0_n_87_12));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r13_reg[11] (.Q(
      execution_unit_0_register_file_0_r13[11]), .QN(), .CK(
      execution_unit_0_register_file_0_n_198), .D(
      execution_unit_0_register_file_0_n_210), .RN(
      execution_unit_0_register_file_0_n_8));
  AND2_X1_LVT execution_unit_0_register_file_0_i_105_246 (.ZN(
      execution_unit_0_register_file_0_n_105_235), .A1(
      execution_unit_0_register_file_0_n_197), .A2(
      execution_unit_0_register_file_0_r13[11]));
  NOR4_X1_LVT execution_unit_0_register_file_0_i_105_247 (.ZN(
      execution_unit_0_register_file_0_n_105_236), .A1(
      execution_unit_0_register_file_0_n_105_224), .A2(
      execution_unit_0_register_file_0_n_105_229), .A3(
      execution_unit_0_register_file_0_n_105_234), .A4(
      execution_unit_0_register_file_0_n_105_235));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_248 (.ZN(
      execution_unit_0_register_file_0_n_105_237), .A1(
      execution_unit_0_register_file_0_n_254), .A2(pc[11]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_101_23 (.ZN(
      execution_unit_0_register_file_0_n_101_12), .A1(
      execution_unit_0_register_file_0_n_101_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[11]), .B1(
      execution_unit_0_register_file_0_r15_wr), .B2(pc_sw[11]));
  INV_X1_LVT execution_unit_0_register_file_0_i_101_24 (.ZN(
      execution_unit_0_register_file_0_n_248), .A(
      execution_unit_0_register_file_0_n_101_12));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r15_reg[11] (.Q(
      execution_unit_0_register_file_0_r15[11]), .QN(), .CK(
      execution_unit_0_register_file_0_n_236), .D(
      execution_unit_0_register_file_0_n_248), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_249 (.ZN(
      execution_unit_0_register_file_0_n_105_238), .A1(
      execution_unit_0_register_file_0_n_235), .A2(
      execution_unit_0_register_file_0_r15[11]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_94_23 (.ZN(
      execution_unit_0_register_file_0_n_94_12), .A1(
      execution_unit_0_register_file_0_n_94_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[11]), .B1(
      execution_unit_0_register_file_0_r14_wr), .B2(pc_sw[11]));
  INV_X1_LVT execution_unit_0_register_file_0_i_94_24 (.ZN(
      execution_unit_0_register_file_0_n_229), .A(
      execution_unit_0_register_file_0_n_94_12));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r14_reg[11] (.Q(
      execution_unit_0_register_file_0_r14[11]), .QN(), .CK(
      execution_unit_0_register_file_0_n_217), .D(
      execution_unit_0_register_file_0_n_229), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_250 (.ZN(
      execution_unit_0_register_file_0_n_105_239), .A1(
      execution_unit_0_register_file_0_n_216), .A2(
      execution_unit_0_register_file_0_r14[11]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_105_251 (.ZN(
      execution_unit_0_reg_src[11]), .A1(
      execution_unit_0_register_file_0_n_105_236), .A2(
      execution_unit_0_register_file_0_n_105_237), .A3(
      execution_unit_0_register_file_0_n_105_238), .A4(
      execution_unit_0_register_file_0_n_105_239));
  HA_X1_LVT execution_unit_0_register_file_0_i_22_11 (.CO(
      execution_unit_0_register_file_0_n_22_11), .S(
      execution_unit_0_register_file_0_reg_incr_val[11]), .A(
      execution_unit_0_reg_src[11]), .B(execution_unit_0_register_file_0_n_22_10));
  HA_X1_LVT execution_unit_0_register_file_0_i_22_12 (.CO(
      execution_unit_0_register_file_0_n_22_12), .S(
      execution_unit_0_register_file_0_reg_incr_val[12]), .A(
      execution_unit_0_reg_src[12]), .B(execution_unit_0_register_file_0_n_22_11));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_24_25 (.ZN(
      execution_unit_0_register_file_0_n_24_13), .A1(
      execution_unit_0_register_file_0_n_24_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[12]), .B1(
      execution_unit_0_register_file_0_r4_wr), .B2(pc_sw[12]));
  INV_X1_LVT execution_unit_0_register_file_0_i_24_26 (.ZN(
      execution_unit_0_register_file_0_n_40), .A(
      execution_unit_0_register_file_0_n_24_13));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r4_reg[12] (.Q(
      execution_unit_0_register_file_0_r4[12]), .QN(), .CK(
      execution_unit_0_register_file_0_n_27), .D(
      execution_unit_0_register_file_0_n_40), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_252 (.ZN(
      execution_unit_0_register_file_0_n_105_240), .A1(
      execution_unit_0_register_file_0_n_24), .A2(
      execution_unit_0_register_file_0_r4[12]));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r3_reg[12] (.Q(
      execution_unit_0_register_file_0_r3[12]), .QN(), .CK(
      execution_unit_0_register_file_0_n_23), .D(pc_sw[12]), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_253 (.ZN(
      execution_unit_0_register_file_0_n_105_241), .A1(
      execution_unit_0_register_file_0_n_22), .A2(
      execution_unit_0_register_file_0_r3[12]));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r2_reg[12] (.Q(
      execution_unit_0_register_file_0_n_3), .QN(), .CK(cpu_mclk), .D(1'b0), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_254 (.ZN(
      execution_unit_0_register_file_0_n_105_242), .A1(
      execution_unit_0_register_file_0_n_21), .A2(
      execution_unit_0_register_file_0_n_3));
  AOI222_X1_LVT execution_unit_0_register_file_0_i_109_22 (.ZN(
      execution_unit_0_register_file_0_n_109_11), .A1(
      execution_unit_0_register_file_0_r1_wr), .A2(pc_sw[12]), .B1(
      execution_unit_0_register_file_0_n_272), .B2(eu_mab[12]), .C1(
      execution_unit_0_register_file_0_n_271), .C2(
      execution_unit_0_register_file_0_n_266));
  INV_X1_LVT execution_unit_0_register_file_0_i_109_23 (.ZN(
      execution_unit_0_register_file_0_n_284), .A(
      execution_unit_0_register_file_0_n_109_11));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r1_reg[12] (.Q(
      execution_unit_0_register_file_0_r1[12]), .QN(), .CK(
      execution_unit_0_register_file_0_n_270), .D(
      execution_unit_0_register_file_0_n_284), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_255 (.ZN(
      execution_unit_0_register_file_0_n_105_243), .A1(
      execution_unit_0_register_file_0_inst_src_in), .A2(
      execution_unit_0_register_file_0_r1[12]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_105_256 (.ZN(
      execution_unit_0_register_file_0_n_105_244), .A1(
      execution_unit_0_register_file_0_n_105_240), .A2(
      execution_unit_0_register_file_0_n_105_241), .A3(
      execution_unit_0_register_file_0_n_105_242), .A4(
      execution_unit_0_register_file_0_n_105_243));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_80_25 (.ZN(
      execution_unit_0_register_file_0_n_80_13), .A1(
      execution_unit_0_register_file_0_n_80_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[12]), .B1(
      execution_unit_0_register_file_0_r12_wr), .B2(pc_sw[12]));
  INV_X1_LVT execution_unit_0_register_file_0_i_80_26 (.ZN(
      execution_unit_0_register_file_0_n_192), .A(
      execution_unit_0_register_file_0_n_80_13));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r12_reg[12] (.Q(
      execution_unit_0_register_file_0_r12[12]), .QN(), .CK(
      execution_unit_0_register_file_0_n_179), .D(
      execution_unit_0_register_file_0_n_192), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_257 (.ZN(
      execution_unit_0_register_file_0_n_105_245), .A1(
      execution_unit_0_register_file_0_n_178), .A2(
      execution_unit_0_register_file_0_r12[12]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_73_25 (.ZN(
      execution_unit_0_register_file_0_n_73_13), .A1(
      execution_unit_0_register_file_0_n_73_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[12]), .B1(
      execution_unit_0_register_file_0_r11_wr), .B2(pc_sw[12]));
  INV_X1_LVT execution_unit_0_register_file_0_i_73_26 (.ZN(
      execution_unit_0_register_file_0_n_173), .A(
      execution_unit_0_register_file_0_n_73_13));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r11_reg[12] (.Q(
      execution_unit_0_register_file_0_r11[12]), .QN(), .CK(
      execution_unit_0_register_file_0_n_160), .D(
      execution_unit_0_register_file_0_n_173), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_258 (.ZN(
      execution_unit_0_register_file_0_n_105_246), .A1(
      execution_unit_0_register_file_0_n_159), .A2(
      execution_unit_0_register_file_0_r11[12]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_66_25 (.ZN(
      execution_unit_0_register_file_0_n_66_13), .A1(
      execution_unit_0_register_file_0_n_66_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[12]), .B1(
      execution_unit_0_register_file_0_r10_wr), .B2(pc_sw[12]));
  INV_X1_LVT execution_unit_0_register_file_0_i_66_26 (.ZN(
      execution_unit_0_register_file_0_n_154), .A(
      execution_unit_0_register_file_0_n_66_13));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r10_reg[12] (.Q(
      execution_unit_0_register_file_0_r10[12]), .QN(), .CK(
      execution_unit_0_register_file_0_n_141), .D(
      execution_unit_0_register_file_0_n_154), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_259 (.ZN(
      execution_unit_0_register_file_0_n_105_247), .A1(
      execution_unit_0_register_file_0_n_140), .A2(
      execution_unit_0_register_file_0_r10[12]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_59_25 (.ZN(
      execution_unit_0_register_file_0_n_59_13), .A1(
      execution_unit_0_register_file_0_n_59_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[12]), .B1(
      execution_unit_0_register_file_0_r9_wr), .B2(pc_sw[12]));
  INV_X1_LVT execution_unit_0_register_file_0_i_59_26 (.ZN(
      execution_unit_0_register_file_0_n_135), .A(
      execution_unit_0_register_file_0_n_59_13));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r9_reg[12] (.Q(
      execution_unit_0_register_file_0_r9[12]), .QN(), .CK(
      execution_unit_0_register_file_0_n_122), .D(
      execution_unit_0_register_file_0_n_135), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_260 (.ZN(
      execution_unit_0_register_file_0_n_105_248), .A1(
      execution_unit_0_register_file_0_n_121), .A2(
      execution_unit_0_register_file_0_r9[12]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_105_261 (.ZN(
      execution_unit_0_register_file_0_n_105_249), .A1(
      execution_unit_0_register_file_0_n_105_245), .A2(
      execution_unit_0_register_file_0_n_105_246), .A3(
      execution_unit_0_register_file_0_n_105_247), .A4(
      execution_unit_0_register_file_0_n_105_248));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_52_25 (.ZN(
      execution_unit_0_register_file_0_n_52_13), .A1(
      execution_unit_0_register_file_0_n_52_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[12]), .B1(
      execution_unit_0_register_file_0_r8_wr), .B2(pc_sw[12]));
  INV_X1_LVT execution_unit_0_register_file_0_i_52_26 (.ZN(
      execution_unit_0_register_file_0_n_116), .A(
      execution_unit_0_register_file_0_n_52_13));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r8_reg[12] (.Q(
      execution_unit_0_register_file_0_r8[12]), .QN(), .CK(
      execution_unit_0_register_file_0_n_103), .D(
      execution_unit_0_register_file_0_n_116), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_262 (.ZN(
      execution_unit_0_register_file_0_n_105_250), .A1(
      execution_unit_0_register_file_0_n_102), .A2(
      execution_unit_0_register_file_0_r8[12]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_45_25 (.ZN(
      execution_unit_0_register_file_0_n_45_13), .A1(
      execution_unit_0_register_file_0_n_45_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[12]), .B1(
      execution_unit_0_register_file_0_r7_wr), .B2(pc_sw[12]));
  INV_X1_LVT execution_unit_0_register_file_0_i_45_26 (.ZN(
      execution_unit_0_register_file_0_n_97), .A(
      execution_unit_0_register_file_0_n_45_13));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r7_reg[12] (.Q(
      execution_unit_0_register_file_0_r7[12]), .QN(), .CK(
      execution_unit_0_register_file_0_n_84), .D(
      execution_unit_0_register_file_0_n_97), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_263 (.ZN(
      execution_unit_0_register_file_0_n_105_251), .A1(
      execution_unit_0_register_file_0_n_83), .A2(
      execution_unit_0_register_file_0_r7[12]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_38_25 (.ZN(
      execution_unit_0_register_file_0_n_38_13), .A1(
      execution_unit_0_register_file_0_n_38_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[12]), .B1(
      execution_unit_0_register_file_0_r6_wr), .B2(pc_sw[12]));
  INV_X1_LVT execution_unit_0_register_file_0_i_38_26 (.ZN(
      execution_unit_0_register_file_0_n_78), .A(
      execution_unit_0_register_file_0_n_38_13));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r6_reg[12] (.Q(
      execution_unit_0_register_file_0_r6[12]), .QN(), .CK(
      execution_unit_0_register_file_0_n_65), .D(
      execution_unit_0_register_file_0_n_78), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_264 (.ZN(
      execution_unit_0_register_file_0_n_105_252), .A1(
      execution_unit_0_register_file_0_n_64), .A2(
      execution_unit_0_register_file_0_r6[12]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_31_25 (.ZN(
      execution_unit_0_register_file_0_n_31_13), .A1(
      execution_unit_0_register_file_0_n_31_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[12]), .B1(
      execution_unit_0_register_file_0_r5_wr), .B2(pc_sw[12]));
  INV_X1_LVT execution_unit_0_register_file_0_i_31_26 (.ZN(
      execution_unit_0_register_file_0_n_59), .A(
      execution_unit_0_register_file_0_n_31_13));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r5_reg[12] (.Q(
      execution_unit_0_register_file_0_r5[12]), .QN(), .CK(
      execution_unit_0_register_file_0_n_46), .D(
      execution_unit_0_register_file_0_n_59), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_265 (.ZN(
      execution_unit_0_register_file_0_n_105_253), .A1(
      execution_unit_0_register_file_0_n_45), .A2(
      execution_unit_0_register_file_0_r5[12]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_105_266 (.ZN(
      execution_unit_0_register_file_0_n_105_254), .A1(
      execution_unit_0_register_file_0_n_105_250), .A2(
      execution_unit_0_register_file_0_n_105_251), .A3(
      execution_unit_0_register_file_0_n_105_252), .A4(
      execution_unit_0_register_file_0_n_105_253));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_87_25 (.ZN(
      execution_unit_0_register_file_0_n_87_13), .A1(
      execution_unit_0_register_file_0_n_87_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[12]), .B1(
      execution_unit_0_register_file_0_r13_wr), .B2(pc_sw[12]));
  INV_X1_LVT execution_unit_0_register_file_0_i_87_26 (.ZN(
      execution_unit_0_register_file_0_n_211), .A(
      execution_unit_0_register_file_0_n_87_13));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r13_reg[12] (.Q(
      execution_unit_0_register_file_0_r13[12]), .QN(), .CK(
      execution_unit_0_register_file_0_n_198), .D(
      execution_unit_0_register_file_0_n_211), .RN(
      execution_unit_0_register_file_0_n_8));
  AND2_X1_LVT execution_unit_0_register_file_0_i_105_267 (.ZN(
      execution_unit_0_register_file_0_n_105_255), .A1(
      execution_unit_0_register_file_0_n_197), .A2(
      execution_unit_0_register_file_0_r13[12]));
  NOR4_X1_LVT execution_unit_0_register_file_0_i_105_268 (.ZN(
      execution_unit_0_register_file_0_n_105_256), .A1(
      execution_unit_0_register_file_0_n_105_244), .A2(
      execution_unit_0_register_file_0_n_105_249), .A3(
      execution_unit_0_register_file_0_n_105_254), .A4(
      execution_unit_0_register_file_0_n_105_255));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_269 (.ZN(
      execution_unit_0_register_file_0_n_105_257), .A1(
      execution_unit_0_register_file_0_n_254), .A2(pc[12]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_101_25 (.ZN(
      execution_unit_0_register_file_0_n_101_13), .A1(
      execution_unit_0_register_file_0_n_101_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[12]), .B1(
      execution_unit_0_register_file_0_r15_wr), .B2(pc_sw[12]));
  INV_X1_LVT execution_unit_0_register_file_0_i_101_26 (.ZN(
      execution_unit_0_register_file_0_n_249), .A(
      execution_unit_0_register_file_0_n_101_13));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r15_reg[12] (.Q(
      execution_unit_0_register_file_0_r15[12]), .QN(), .CK(
      execution_unit_0_register_file_0_n_236), .D(
      execution_unit_0_register_file_0_n_249), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_270 (.ZN(
      execution_unit_0_register_file_0_n_105_258), .A1(
      execution_unit_0_register_file_0_n_235), .A2(
      execution_unit_0_register_file_0_r15[12]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_94_25 (.ZN(
      execution_unit_0_register_file_0_n_94_13), .A1(
      execution_unit_0_register_file_0_n_94_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[12]), .B1(
      execution_unit_0_register_file_0_r14_wr), .B2(pc_sw[12]));
  INV_X1_LVT execution_unit_0_register_file_0_i_94_26 (.ZN(
      execution_unit_0_register_file_0_n_230), .A(
      execution_unit_0_register_file_0_n_94_13));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r14_reg[12] (.Q(
      execution_unit_0_register_file_0_r14[12]), .QN(), .CK(
      execution_unit_0_register_file_0_n_217), .D(
      execution_unit_0_register_file_0_n_230), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_271 (.ZN(
      execution_unit_0_register_file_0_n_105_259), .A1(
      execution_unit_0_register_file_0_n_216), .A2(
      execution_unit_0_register_file_0_r14[12]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_105_272 (.ZN(
      execution_unit_0_reg_src[12]), .A1(
      execution_unit_0_register_file_0_n_105_256), .A2(
      execution_unit_0_register_file_0_n_105_257), .A3(
      execution_unit_0_register_file_0_n_105_258), .A4(
      execution_unit_0_register_file_0_n_105_259));
  HA_X1_LVT execution_unit_0_register_file_0_i_106_11 (.CO(
      execution_unit_0_register_file_0_n_106_10), .S(
      execution_unit_0_register_file_0_n_266), .A(execution_unit_0_reg_src[12]), 
      .B(execution_unit_0_register_file_0_n_106_9));
  HA_X1_LVT execution_unit_0_register_file_0_i_106_12 (.CO(
      execution_unit_0_register_file_0_n_106_11), .S(
      execution_unit_0_register_file_0_n_267), .A(execution_unit_0_reg_src[13]), 
      .B(execution_unit_0_register_file_0_n_106_10));
  AOI222_X1_LVT execution_unit_0_register_file_0_i_109_24 (.ZN(
      execution_unit_0_register_file_0_n_109_12), .A1(
      execution_unit_0_register_file_0_r1_wr), .A2(pc_sw[13]), .B1(
      execution_unit_0_register_file_0_n_272), .B2(eu_mab[13]), .C1(
      execution_unit_0_register_file_0_n_271), .C2(
      execution_unit_0_register_file_0_n_267));
  INV_X1_LVT execution_unit_0_register_file_0_i_109_25 (.ZN(
      execution_unit_0_register_file_0_n_285), .A(
      execution_unit_0_register_file_0_n_109_12));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r1_reg[13] (.Q(
      execution_unit_0_register_file_0_r1[13]), .QN(), .CK(
      execution_unit_0_register_file_0_n_270), .D(
      execution_unit_0_register_file_0_n_285), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_276 (.ZN(
      execution_unit_0_register_file_0_n_105_263), .A1(
      execution_unit_0_register_file_0_inst_src_in), .A2(
      execution_unit_0_register_file_0_r1[13]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_105_277 (.ZN(
      execution_unit_0_register_file_0_n_105_264), .A1(
      execution_unit_0_register_file_0_n_105_260), .A2(
      execution_unit_0_register_file_0_n_105_261), .A3(
      execution_unit_0_register_file_0_n_105_262), .A4(
      execution_unit_0_register_file_0_n_105_263));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_80_27 (.ZN(
      execution_unit_0_register_file_0_n_80_14), .A1(
      execution_unit_0_register_file_0_n_80_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[13]), .B1(
      execution_unit_0_register_file_0_r12_wr), .B2(pc_sw[13]));
  INV_X1_LVT execution_unit_0_register_file_0_i_80_28 (.ZN(
      execution_unit_0_register_file_0_n_193), .A(
      execution_unit_0_register_file_0_n_80_14));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r12_reg[13] (.Q(
      execution_unit_0_register_file_0_r12[13]), .QN(), .CK(
      execution_unit_0_register_file_0_n_179), .D(
      execution_unit_0_register_file_0_n_193), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_278 (.ZN(
      execution_unit_0_register_file_0_n_105_265), .A1(
      execution_unit_0_register_file_0_n_178), .A2(
      execution_unit_0_register_file_0_r12[13]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_73_27 (.ZN(
      execution_unit_0_register_file_0_n_73_14), .A1(
      execution_unit_0_register_file_0_n_73_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[13]), .B1(
      execution_unit_0_register_file_0_r11_wr), .B2(pc_sw[13]));
  INV_X1_LVT execution_unit_0_register_file_0_i_73_28 (.ZN(
      execution_unit_0_register_file_0_n_174), .A(
      execution_unit_0_register_file_0_n_73_14));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r11_reg[13] (.Q(
      execution_unit_0_register_file_0_r11[13]), .QN(), .CK(
      execution_unit_0_register_file_0_n_160), .D(
      execution_unit_0_register_file_0_n_174), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_279 (.ZN(
      execution_unit_0_register_file_0_n_105_266), .A1(
      execution_unit_0_register_file_0_n_159), .A2(
      execution_unit_0_register_file_0_r11[13]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_66_27 (.ZN(
      execution_unit_0_register_file_0_n_66_14), .A1(
      execution_unit_0_register_file_0_n_66_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[13]), .B1(
      execution_unit_0_register_file_0_r10_wr), .B2(pc_sw[13]));
  INV_X1_LVT execution_unit_0_register_file_0_i_66_28 (.ZN(
      execution_unit_0_register_file_0_n_155), .A(
      execution_unit_0_register_file_0_n_66_14));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r10_reg[13] (.Q(
      execution_unit_0_register_file_0_r10[13]), .QN(), .CK(
      execution_unit_0_register_file_0_n_141), .D(
      execution_unit_0_register_file_0_n_155), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_280 (.ZN(
      execution_unit_0_register_file_0_n_105_267), .A1(
      execution_unit_0_register_file_0_n_140), .A2(
      execution_unit_0_register_file_0_r10[13]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_59_27 (.ZN(
      execution_unit_0_register_file_0_n_59_14), .A1(
      execution_unit_0_register_file_0_n_59_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[13]), .B1(
      execution_unit_0_register_file_0_r9_wr), .B2(pc_sw[13]));
  INV_X1_LVT execution_unit_0_register_file_0_i_59_28 (.ZN(
      execution_unit_0_register_file_0_n_136), .A(
      execution_unit_0_register_file_0_n_59_14));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r9_reg[13] (.Q(
      execution_unit_0_register_file_0_r9[13]), .QN(), .CK(
      execution_unit_0_register_file_0_n_122), .D(
      execution_unit_0_register_file_0_n_136), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_281 (.ZN(
      execution_unit_0_register_file_0_n_105_268), .A1(
      execution_unit_0_register_file_0_n_121), .A2(
      execution_unit_0_register_file_0_r9[13]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_105_282 (.ZN(
      execution_unit_0_register_file_0_n_105_269), .A1(
      execution_unit_0_register_file_0_n_105_265), .A2(
      execution_unit_0_register_file_0_n_105_266), .A3(
      execution_unit_0_register_file_0_n_105_267), .A4(
      execution_unit_0_register_file_0_n_105_268));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_52_27 (.ZN(
      execution_unit_0_register_file_0_n_52_14), .A1(
      execution_unit_0_register_file_0_n_52_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[13]), .B1(
      execution_unit_0_register_file_0_r8_wr), .B2(pc_sw[13]));
  INV_X1_LVT execution_unit_0_register_file_0_i_52_28 (.ZN(
      execution_unit_0_register_file_0_n_117), .A(
      execution_unit_0_register_file_0_n_52_14));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r8_reg[13] (.Q(
      execution_unit_0_register_file_0_r8[13]), .QN(), .CK(
      execution_unit_0_register_file_0_n_103), .D(
      execution_unit_0_register_file_0_n_117), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_283 (.ZN(
      execution_unit_0_register_file_0_n_105_270), .A1(
      execution_unit_0_register_file_0_n_102), .A2(
      execution_unit_0_register_file_0_r8[13]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_45_27 (.ZN(
      execution_unit_0_register_file_0_n_45_14), .A1(
      execution_unit_0_register_file_0_n_45_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[13]), .B1(
      execution_unit_0_register_file_0_r7_wr), .B2(pc_sw[13]));
  INV_X1_LVT execution_unit_0_register_file_0_i_45_28 (.ZN(
      execution_unit_0_register_file_0_n_98), .A(
      execution_unit_0_register_file_0_n_45_14));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r7_reg[13] (.Q(
      execution_unit_0_register_file_0_r7[13]), .QN(), .CK(
      execution_unit_0_register_file_0_n_84), .D(
      execution_unit_0_register_file_0_n_98), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_284 (.ZN(
      execution_unit_0_register_file_0_n_105_271), .A1(
      execution_unit_0_register_file_0_n_83), .A2(
      execution_unit_0_register_file_0_r7[13]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_38_27 (.ZN(
      execution_unit_0_register_file_0_n_38_14), .A1(
      execution_unit_0_register_file_0_n_38_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[13]), .B1(
      execution_unit_0_register_file_0_r6_wr), .B2(pc_sw[13]));
  INV_X1_LVT execution_unit_0_register_file_0_i_38_28 (.ZN(
      execution_unit_0_register_file_0_n_79), .A(
      execution_unit_0_register_file_0_n_38_14));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r6_reg[13] (.Q(
      execution_unit_0_register_file_0_r6[13]), .QN(), .CK(
      execution_unit_0_register_file_0_n_65), .D(
      execution_unit_0_register_file_0_n_79), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_285 (.ZN(
      execution_unit_0_register_file_0_n_105_272), .A1(
      execution_unit_0_register_file_0_n_64), .A2(
      execution_unit_0_register_file_0_r6[13]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_31_27 (.ZN(
      execution_unit_0_register_file_0_n_31_14), .A1(
      execution_unit_0_register_file_0_n_31_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[13]), .B1(
      execution_unit_0_register_file_0_r5_wr), .B2(pc_sw[13]));
  INV_X1_LVT execution_unit_0_register_file_0_i_31_28 (.ZN(
      execution_unit_0_register_file_0_n_60), .A(
      execution_unit_0_register_file_0_n_31_14));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r5_reg[13] (.Q(
      execution_unit_0_register_file_0_r5[13]), .QN(), .CK(
      execution_unit_0_register_file_0_n_46), .D(
      execution_unit_0_register_file_0_n_60), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_286 (.ZN(
      execution_unit_0_register_file_0_n_105_273), .A1(
      execution_unit_0_register_file_0_n_45), .A2(
      execution_unit_0_register_file_0_r5[13]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_105_287 (.ZN(
      execution_unit_0_register_file_0_n_105_274), .A1(
      execution_unit_0_register_file_0_n_105_270), .A2(
      execution_unit_0_register_file_0_n_105_271), .A3(
      execution_unit_0_register_file_0_n_105_272), .A4(
      execution_unit_0_register_file_0_n_105_273));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_87_27 (.ZN(
      execution_unit_0_register_file_0_n_87_14), .A1(
      execution_unit_0_register_file_0_n_87_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[13]), .B1(
      execution_unit_0_register_file_0_r13_wr), .B2(pc_sw[13]));
  INV_X1_LVT execution_unit_0_register_file_0_i_87_28 (.ZN(
      execution_unit_0_register_file_0_n_212), .A(
      execution_unit_0_register_file_0_n_87_14));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r13_reg[13] (.Q(
      execution_unit_0_register_file_0_r13[13]), .QN(), .CK(
      execution_unit_0_register_file_0_n_198), .D(
      execution_unit_0_register_file_0_n_212), .RN(
      execution_unit_0_register_file_0_n_8));
  AND2_X1_LVT execution_unit_0_register_file_0_i_105_288 (.ZN(
      execution_unit_0_register_file_0_n_105_275), .A1(
      execution_unit_0_register_file_0_n_197), .A2(
      execution_unit_0_register_file_0_r13[13]));
  NOR4_X1_LVT execution_unit_0_register_file_0_i_105_289 (.ZN(
      execution_unit_0_register_file_0_n_105_276), .A1(
      execution_unit_0_register_file_0_n_105_264), .A2(
      execution_unit_0_register_file_0_n_105_269), .A3(
      execution_unit_0_register_file_0_n_105_274), .A4(
      execution_unit_0_register_file_0_n_105_275));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_290 (.ZN(
      execution_unit_0_register_file_0_n_105_277), .A1(
      execution_unit_0_register_file_0_n_254), .A2(pc[13]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_101_27 (.ZN(
      execution_unit_0_register_file_0_n_101_14), .A1(
      execution_unit_0_register_file_0_n_101_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[13]), .B1(
      execution_unit_0_register_file_0_r15_wr), .B2(pc_sw[13]));
  INV_X1_LVT execution_unit_0_register_file_0_i_101_28 (.ZN(
      execution_unit_0_register_file_0_n_250), .A(
      execution_unit_0_register_file_0_n_101_14));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r15_reg[13] (.Q(
      execution_unit_0_register_file_0_r15[13]), .QN(), .CK(
      execution_unit_0_register_file_0_n_236), .D(
      execution_unit_0_register_file_0_n_250), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_291 (.ZN(
      execution_unit_0_register_file_0_n_105_278), .A1(
      execution_unit_0_register_file_0_n_235), .A2(
      execution_unit_0_register_file_0_r15[13]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_94_27 (.ZN(
      execution_unit_0_register_file_0_n_94_14), .A1(
      execution_unit_0_register_file_0_n_94_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[13]), .B1(
      execution_unit_0_register_file_0_r14_wr), .B2(pc_sw[13]));
  INV_X1_LVT execution_unit_0_register_file_0_i_94_28 (.ZN(
      execution_unit_0_register_file_0_n_231), .A(
      execution_unit_0_register_file_0_n_94_14));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r14_reg[13] (.Q(
      execution_unit_0_register_file_0_r14[13]), .QN(), .CK(
      execution_unit_0_register_file_0_n_217), .D(
      execution_unit_0_register_file_0_n_231), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_292 (.ZN(
      execution_unit_0_register_file_0_n_105_279), .A1(
      execution_unit_0_register_file_0_n_216), .A2(
      execution_unit_0_register_file_0_r14[13]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_105_293 (.ZN(
      execution_unit_0_reg_src[13]), .A1(
      execution_unit_0_register_file_0_n_105_276), .A2(
      execution_unit_0_register_file_0_n_105_277), .A3(
      execution_unit_0_register_file_0_n_105_278), .A4(
      execution_unit_0_register_file_0_n_105_279));
  HA_X1_LVT execution_unit_0_register_file_0_i_22_13 (.CO(
      execution_unit_0_register_file_0_n_22_13), .S(
      execution_unit_0_register_file_0_reg_incr_val[13]), .A(
      execution_unit_0_reg_src[13]), .B(execution_unit_0_register_file_0_n_22_12));
  HA_X1_LVT execution_unit_0_register_file_0_i_22_14 (.CO(
      execution_unit_0_register_file_0_n_22_14), .S(
      execution_unit_0_register_file_0_reg_incr_val[14]), .A(
      execution_unit_0_reg_src[14]), .B(execution_unit_0_register_file_0_n_22_13));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_24_29 (.ZN(
      execution_unit_0_register_file_0_n_24_15), .A1(
      execution_unit_0_register_file_0_n_24_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[14]), .B1(
      execution_unit_0_register_file_0_r4_wr), .B2(pc_sw[14]));
  INV_X1_LVT execution_unit_0_register_file_0_i_24_30 (.ZN(
      execution_unit_0_register_file_0_n_42), .A(
      execution_unit_0_register_file_0_n_24_15));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r4_reg[14] (.Q(
      execution_unit_0_register_file_0_r4[14]), .QN(), .CK(
      execution_unit_0_register_file_0_n_27), .D(
      execution_unit_0_register_file_0_n_42), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_294 (.ZN(
      execution_unit_0_register_file_0_n_105_280), .A1(
      execution_unit_0_register_file_0_n_24), .A2(
      execution_unit_0_register_file_0_r4[14]));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r3_reg[14] (.Q(
      execution_unit_0_register_file_0_r3[14]), .QN(), .CK(
      execution_unit_0_register_file_0_n_23), .D(pc_sw[14]), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_295 (.ZN(
      execution_unit_0_register_file_0_n_105_281), .A1(
      execution_unit_0_register_file_0_n_22), .A2(
      execution_unit_0_register_file_0_r3[14]));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r2_reg[14] (.Q(
      execution_unit_0_register_file_0_n_1), .QN(), .CK(cpu_mclk), .D(1'b0), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_296 (.ZN(
      execution_unit_0_register_file_0_n_105_282), .A1(
      execution_unit_0_register_file_0_n_21), .A2(
      execution_unit_0_register_file_0_n_1));
  AOI222_X1_LVT execution_unit_0_register_file_0_i_109_26 (.ZN(
      execution_unit_0_register_file_0_n_109_13), .A1(
      execution_unit_0_register_file_0_r1_wr), .A2(pc_sw[14]), .B1(
      execution_unit_0_register_file_0_n_272), .B2(eu_mab[14]), .C1(
      execution_unit_0_register_file_0_n_271), .C2(
      execution_unit_0_register_file_0_n_268));
  INV_X1_LVT execution_unit_0_register_file_0_i_109_27 (.ZN(
      execution_unit_0_register_file_0_n_286), .A(
      execution_unit_0_register_file_0_n_109_13));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r1_reg[14] (.Q(
      execution_unit_0_register_file_0_r1[14]), .QN(), .CK(
      execution_unit_0_register_file_0_n_270), .D(
      execution_unit_0_register_file_0_n_286), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_297 (.ZN(
      execution_unit_0_register_file_0_n_105_283), .A1(
      execution_unit_0_register_file_0_inst_src_in), .A2(
      execution_unit_0_register_file_0_r1[14]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_105_298 (.ZN(
      execution_unit_0_register_file_0_n_105_284), .A1(
      execution_unit_0_register_file_0_n_105_280), .A2(
      execution_unit_0_register_file_0_n_105_281), .A3(
      execution_unit_0_register_file_0_n_105_282), .A4(
      execution_unit_0_register_file_0_n_105_283));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_80_29 (.ZN(
      execution_unit_0_register_file_0_n_80_15), .A1(
      execution_unit_0_register_file_0_n_80_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[14]), .B1(
      execution_unit_0_register_file_0_r12_wr), .B2(pc_sw[14]));
  INV_X1_LVT execution_unit_0_register_file_0_i_80_30 (.ZN(
      execution_unit_0_register_file_0_n_194), .A(
      execution_unit_0_register_file_0_n_80_15));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r12_reg[14] (.Q(
      execution_unit_0_register_file_0_r12[14]), .QN(), .CK(
      execution_unit_0_register_file_0_n_179), .D(
      execution_unit_0_register_file_0_n_194), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_299 (.ZN(
      execution_unit_0_register_file_0_n_105_285), .A1(
      execution_unit_0_register_file_0_n_178), .A2(
      execution_unit_0_register_file_0_r12[14]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_73_29 (.ZN(
      execution_unit_0_register_file_0_n_73_15), .A1(
      execution_unit_0_register_file_0_n_73_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[14]), .B1(
      execution_unit_0_register_file_0_r11_wr), .B2(pc_sw[14]));
  INV_X1_LVT execution_unit_0_register_file_0_i_73_30 (.ZN(
      execution_unit_0_register_file_0_n_175), .A(
      execution_unit_0_register_file_0_n_73_15));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r11_reg[14] (.Q(
      execution_unit_0_register_file_0_r11[14]), .QN(), .CK(
      execution_unit_0_register_file_0_n_160), .D(
      execution_unit_0_register_file_0_n_175), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_300 (.ZN(
      execution_unit_0_register_file_0_n_105_286), .A1(
      execution_unit_0_register_file_0_n_159), .A2(
      execution_unit_0_register_file_0_r11[14]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_66_29 (.ZN(
      execution_unit_0_register_file_0_n_66_15), .A1(
      execution_unit_0_register_file_0_n_66_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[14]), .B1(
      execution_unit_0_register_file_0_r10_wr), .B2(pc_sw[14]));
  INV_X1_LVT execution_unit_0_register_file_0_i_66_30 (.ZN(
      execution_unit_0_register_file_0_n_156), .A(
      execution_unit_0_register_file_0_n_66_15));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r10_reg[14] (.Q(
      execution_unit_0_register_file_0_r10[14]), .QN(), .CK(
      execution_unit_0_register_file_0_n_141), .D(
      execution_unit_0_register_file_0_n_156), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_301 (.ZN(
      execution_unit_0_register_file_0_n_105_287), .A1(
      execution_unit_0_register_file_0_n_140), .A2(
      execution_unit_0_register_file_0_r10[14]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_59_29 (.ZN(
      execution_unit_0_register_file_0_n_59_15), .A1(
      execution_unit_0_register_file_0_n_59_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[14]), .B1(
      execution_unit_0_register_file_0_r9_wr), .B2(pc_sw[14]));
  INV_X1_LVT execution_unit_0_register_file_0_i_59_30 (.ZN(
      execution_unit_0_register_file_0_n_137), .A(
      execution_unit_0_register_file_0_n_59_15));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r9_reg[14] (.Q(
      execution_unit_0_register_file_0_r9[14]), .QN(), .CK(
      execution_unit_0_register_file_0_n_122), .D(
      execution_unit_0_register_file_0_n_137), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_302 (.ZN(
      execution_unit_0_register_file_0_n_105_288), .A1(
      execution_unit_0_register_file_0_n_121), .A2(
      execution_unit_0_register_file_0_r9[14]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_105_303 (.ZN(
      execution_unit_0_register_file_0_n_105_289), .A1(
      execution_unit_0_register_file_0_n_105_285), .A2(
      execution_unit_0_register_file_0_n_105_286), .A3(
      execution_unit_0_register_file_0_n_105_287), .A4(
      execution_unit_0_register_file_0_n_105_288));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_52_29 (.ZN(
      execution_unit_0_register_file_0_n_52_15), .A1(
      execution_unit_0_register_file_0_n_52_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[14]), .B1(
      execution_unit_0_register_file_0_r8_wr), .B2(pc_sw[14]));
  INV_X1_LVT execution_unit_0_register_file_0_i_52_30 (.ZN(
      execution_unit_0_register_file_0_n_118), .A(
      execution_unit_0_register_file_0_n_52_15));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r8_reg[14] (.Q(
      execution_unit_0_register_file_0_r8[14]), .QN(), .CK(
      execution_unit_0_register_file_0_n_103), .D(
      execution_unit_0_register_file_0_n_118), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_304 (.ZN(
      execution_unit_0_register_file_0_n_105_290), .A1(
      execution_unit_0_register_file_0_n_102), .A2(
      execution_unit_0_register_file_0_r8[14]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_45_29 (.ZN(
      execution_unit_0_register_file_0_n_45_15), .A1(
      execution_unit_0_register_file_0_n_45_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[14]), .B1(
      execution_unit_0_register_file_0_r7_wr), .B2(pc_sw[14]));
  INV_X1_LVT execution_unit_0_register_file_0_i_45_30 (.ZN(
      execution_unit_0_register_file_0_n_99), .A(
      execution_unit_0_register_file_0_n_45_15));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r7_reg[14] (.Q(
      execution_unit_0_register_file_0_r7[14]), .QN(), .CK(
      execution_unit_0_register_file_0_n_84), .D(
      execution_unit_0_register_file_0_n_99), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_305 (.ZN(
      execution_unit_0_register_file_0_n_105_291), .A1(
      execution_unit_0_register_file_0_n_83), .A2(
      execution_unit_0_register_file_0_r7[14]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_38_29 (.ZN(
      execution_unit_0_register_file_0_n_38_15), .A1(
      execution_unit_0_register_file_0_n_38_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[14]), .B1(
      execution_unit_0_register_file_0_r6_wr), .B2(pc_sw[14]));
  INV_X1_LVT execution_unit_0_register_file_0_i_38_30 (.ZN(
      execution_unit_0_register_file_0_n_80), .A(
      execution_unit_0_register_file_0_n_38_15));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r6_reg[14] (.Q(
      execution_unit_0_register_file_0_r6[14]), .QN(), .CK(
      execution_unit_0_register_file_0_n_65), .D(
      execution_unit_0_register_file_0_n_80), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_306 (.ZN(
      execution_unit_0_register_file_0_n_105_292), .A1(
      execution_unit_0_register_file_0_n_64), .A2(
      execution_unit_0_register_file_0_r6[14]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_31_29 (.ZN(
      execution_unit_0_register_file_0_n_31_15), .A1(
      execution_unit_0_register_file_0_n_31_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[14]), .B1(
      execution_unit_0_register_file_0_r5_wr), .B2(pc_sw[14]));
  INV_X1_LVT execution_unit_0_register_file_0_i_31_30 (.ZN(
      execution_unit_0_register_file_0_n_61), .A(
      execution_unit_0_register_file_0_n_31_15));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r5_reg[14] (.Q(
      execution_unit_0_register_file_0_r5[14]), .QN(), .CK(
      execution_unit_0_register_file_0_n_46), .D(
      execution_unit_0_register_file_0_n_61), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_307 (.ZN(
      execution_unit_0_register_file_0_n_105_293), .A1(
      execution_unit_0_register_file_0_n_45), .A2(
      execution_unit_0_register_file_0_r5[14]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_105_308 (.ZN(
      execution_unit_0_register_file_0_n_105_294), .A1(
      execution_unit_0_register_file_0_n_105_290), .A2(
      execution_unit_0_register_file_0_n_105_291), .A3(
      execution_unit_0_register_file_0_n_105_292), .A4(
      execution_unit_0_register_file_0_n_105_293));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_87_29 (.ZN(
      execution_unit_0_register_file_0_n_87_15), .A1(
      execution_unit_0_register_file_0_n_87_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[14]), .B1(
      execution_unit_0_register_file_0_r13_wr), .B2(pc_sw[14]));
  INV_X1_LVT execution_unit_0_register_file_0_i_87_30 (.ZN(
      execution_unit_0_register_file_0_n_213), .A(
      execution_unit_0_register_file_0_n_87_15));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r13_reg[14] (.Q(
      execution_unit_0_register_file_0_r13[14]), .QN(), .CK(
      execution_unit_0_register_file_0_n_198), .D(
      execution_unit_0_register_file_0_n_213), .RN(
      execution_unit_0_register_file_0_n_8));
  AND2_X1_LVT execution_unit_0_register_file_0_i_105_309 (.ZN(
      execution_unit_0_register_file_0_n_105_295), .A1(
      execution_unit_0_register_file_0_n_197), .A2(
      execution_unit_0_register_file_0_r13[14]));
  NOR4_X1_LVT execution_unit_0_register_file_0_i_105_310 (.ZN(
      execution_unit_0_register_file_0_n_105_296), .A1(
      execution_unit_0_register_file_0_n_105_284), .A2(
      execution_unit_0_register_file_0_n_105_289), .A3(
      execution_unit_0_register_file_0_n_105_294), .A4(
      execution_unit_0_register_file_0_n_105_295));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_311 (.ZN(
      execution_unit_0_register_file_0_n_105_297), .A1(
      execution_unit_0_register_file_0_n_254), .A2(pc[14]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_101_29 (.ZN(
      execution_unit_0_register_file_0_n_101_15), .A1(
      execution_unit_0_register_file_0_n_101_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[14]), .B1(
      execution_unit_0_register_file_0_r15_wr), .B2(pc_sw[14]));
  INV_X1_LVT execution_unit_0_register_file_0_i_101_30 (.ZN(
      execution_unit_0_register_file_0_n_251), .A(
      execution_unit_0_register_file_0_n_101_15));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r15_reg[14] (.Q(
      execution_unit_0_register_file_0_r15[14]), .QN(), .CK(
      execution_unit_0_register_file_0_n_236), .D(
      execution_unit_0_register_file_0_n_251), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_312 (.ZN(
      execution_unit_0_register_file_0_n_105_298), .A1(
      execution_unit_0_register_file_0_n_235), .A2(
      execution_unit_0_register_file_0_r15[14]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_94_29 (.ZN(
      execution_unit_0_register_file_0_n_94_15), .A1(
      execution_unit_0_register_file_0_n_94_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[14]), .B1(
      execution_unit_0_register_file_0_r14_wr), .B2(pc_sw[14]));
  INV_X1_LVT execution_unit_0_register_file_0_i_94_30 (.ZN(
      execution_unit_0_register_file_0_n_232), .A(
      execution_unit_0_register_file_0_n_94_15));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r14_reg[14] (.Q(
      execution_unit_0_register_file_0_r14[14]), .QN(), .CK(
      execution_unit_0_register_file_0_n_217), .D(
      execution_unit_0_register_file_0_n_232), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_313 (.ZN(
      execution_unit_0_register_file_0_n_105_299), .A1(
      execution_unit_0_register_file_0_n_216), .A2(
      execution_unit_0_register_file_0_r14[14]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_105_314 (.ZN(
      execution_unit_0_reg_src[14]), .A1(
      execution_unit_0_register_file_0_n_105_296), .A2(
      execution_unit_0_register_file_0_n_105_297), .A3(
      execution_unit_0_register_file_0_n_105_298), .A4(
      execution_unit_0_register_file_0_n_105_299));
  HA_X1_LVT execution_unit_0_register_file_0_i_106_13 (.CO(
      execution_unit_0_register_file_0_n_106_12), .S(
      execution_unit_0_register_file_0_n_268), .A(execution_unit_0_reg_src[14]), 
      .B(execution_unit_0_register_file_0_n_106_11));
  XNOR2_X1_LVT execution_unit_0_register_file_0_i_106_14 (.ZN(
      execution_unit_0_register_file_0_n_106_13), .A(
      execution_unit_0_reg_src[15]), .B(
      execution_unit_0_register_file_0_n_106_12));
  INV_X1_LVT execution_unit_0_register_file_0_i_106_15 (.ZN(
      execution_unit_0_register_file_0_n_269), .A(
      execution_unit_0_register_file_0_n_106_13));
  AOI222_X1_LVT execution_unit_0_register_file_0_i_109_28 (.ZN(
      execution_unit_0_register_file_0_n_109_14), .A1(
      execution_unit_0_register_file_0_r1_wr), .A2(pc_sw[15]), .B1(
      execution_unit_0_register_file_0_n_272), .B2(eu_mab[15]), .C1(
      execution_unit_0_register_file_0_n_271), .C2(
      execution_unit_0_register_file_0_n_269));
  INV_X1_LVT execution_unit_0_register_file_0_i_109_29 (.ZN(
      execution_unit_0_register_file_0_n_287), .A(
      execution_unit_0_register_file_0_n_109_14));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r1_reg[15] (.Q(
      execution_unit_0_register_file_0_r1[15]), .QN(), .CK(
      execution_unit_0_register_file_0_n_270), .D(
      execution_unit_0_register_file_0_n_287), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_318 (.ZN(
      execution_unit_0_register_file_0_n_105_303), .A1(
      execution_unit_0_register_file_0_inst_src_in), .A2(
      execution_unit_0_register_file_0_r1[15]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_105_319 (.ZN(
      execution_unit_0_register_file_0_n_105_304), .A1(
      execution_unit_0_register_file_0_n_105_300), .A2(
      execution_unit_0_register_file_0_n_105_301), .A3(
      execution_unit_0_register_file_0_n_105_302), .A4(
      execution_unit_0_register_file_0_n_105_303));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_80_31 (.ZN(
      execution_unit_0_register_file_0_n_80_16), .A1(
      execution_unit_0_register_file_0_n_80_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[15]), .B1(
      execution_unit_0_register_file_0_r12_wr), .B2(pc_sw[15]));
  INV_X1_LVT execution_unit_0_register_file_0_i_80_32 (.ZN(
      execution_unit_0_register_file_0_n_195), .A(
      execution_unit_0_register_file_0_n_80_16));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r12_reg[15] (.Q(
      execution_unit_0_register_file_0_r12[15]), .QN(), .CK(
      execution_unit_0_register_file_0_n_179), .D(
      execution_unit_0_register_file_0_n_195), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_320 (.ZN(
      execution_unit_0_register_file_0_n_105_305), .A1(
      execution_unit_0_register_file_0_n_178), .A2(
      execution_unit_0_register_file_0_r12[15]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_73_31 (.ZN(
      execution_unit_0_register_file_0_n_73_16), .A1(
      execution_unit_0_register_file_0_n_73_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[15]), .B1(
      execution_unit_0_register_file_0_r11_wr), .B2(pc_sw[15]));
  INV_X1_LVT execution_unit_0_register_file_0_i_73_32 (.ZN(
      execution_unit_0_register_file_0_n_176), .A(
      execution_unit_0_register_file_0_n_73_16));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r11_reg[15] (.Q(
      execution_unit_0_register_file_0_r11[15]), .QN(), .CK(
      execution_unit_0_register_file_0_n_160), .D(
      execution_unit_0_register_file_0_n_176), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_321 (.ZN(
      execution_unit_0_register_file_0_n_105_306), .A1(
      execution_unit_0_register_file_0_n_159), .A2(
      execution_unit_0_register_file_0_r11[15]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_66_31 (.ZN(
      execution_unit_0_register_file_0_n_66_16), .A1(
      execution_unit_0_register_file_0_n_66_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[15]), .B1(
      execution_unit_0_register_file_0_r10_wr), .B2(pc_sw[15]));
  INV_X1_LVT execution_unit_0_register_file_0_i_66_32 (.ZN(
      execution_unit_0_register_file_0_n_157), .A(
      execution_unit_0_register_file_0_n_66_16));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r10_reg[15] (.Q(
      execution_unit_0_register_file_0_r10[15]), .QN(), .CK(
      execution_unit_0_register_file_0_n_141), .D(
      execution_unit_0_register_file_0_n_157), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_322 (.ZN(
      execution_unit_0_register_file_0_n_105_307), .A1(
      execution_unit_0_register_file_0_n_140), .A2(
      execution_unit_0_register_file_0_r10[15]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_59_31 (.ZN(
      execution_unit_0_register_file_0_n_59_16), .A1(
      execution_unit_0_register_file_0_n_59_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[15]), .B1(
      execution_unit_0_register_file_0_r9_wr), .B2(pc_sw[15]));
  INV_X1_LVT execution_unit_0_register_file_0_i_59_32 (.ZN(
      execution_unit_0_register_file_0_n_138), .A(
      execution_unit_0_register_file_0_n_59_16));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r9_reg[15] (.Q(
      execution_unit_0_register_file_0_r9[15]), .QN(), .CK(
      execution_unit_0_register_file_0_n_122), .D(
      execution_unit_0_register_file_0_n_138), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_323 (.ZN(
      execution_unit_0_register_file_0_n_105_308), .A1(
      execution_unit_0_register_file_0_n_121), .A2(
      execution_unit_0_register_file_0_r9[15]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_105_324 (.ZN(
      execution_unit_0_register_file_0_n_105_309), .A1(
      execution_unit_0_register_file_0_n_105_305), .A2(
      execution_unit_0_register_file_0_n_105_306), .A3(
      execution_unit_0_register_file_0_n_105_307), .A4(
      execution_unit_0_register_file_0_n_105_308));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_52_31 (.ZN(
      execution_unit_0_register_file_0_n_52_16), .A1(
      execution_unit_0_register_file_0_n_52_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[15]), .B1(
      execution_unit_0_register_file_0_r8_wr), .B2(pc_sw[15]));
  INV_X1_LVT execution_unit_0_register_file_0_i_52_32 (.ZN(
      execution_unit_0_register_file_0_n_119), .A(
      execution_unit_0_register_file_0_n_52_16));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r8_reg[15] (.Q(
      execution_unit_0_register_file_0_r8[15]), .QN(), .CK(
      execution_unit_0_register_file_0_n_103), .D(
      execution_unit_0_register_file_0_n_119), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_325 (.ZN(
      execution_unit_0_register_file_0_n_105_310), .A1(
      execution_unit_0_register_file_0_n_102), .A2(
      execution_unit_0_register_file_0_r8[15]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_45_31 (.ZN(
      execution_unit_0_register_file_0_n_45_16), .A1(
      execution_unit_0_register_file_0_n_45_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[15]), .B1(
      execution_unit_0_register_file_0_r7_wr), .B2(pc_sw[15]));
  INV_X1_LVT execution_unit_0_register_file_0_i_45_32 (.ZN(
      execution_unit_0_register_file_0_n_100), .A(
      execution_unit_0_register_file_0_n_45_16));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r7_reg[15] (.Q(
      execution_unit_0_register_file_0_r7[15]), .QN(), .CK(
      execution_unit_0_register_file_0_n_84), .D(
      execution_unit_0_register_file_0_n_100), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_326 (.ZN(
      execution_unit_0_register_file_0_n_105_311), .A1(
      execution_unit_0_register_file_0_n_83), .A2(
      execution_unit_0_register_file_0_r7[15]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_38_31 (.ZN(
      execution_unit_0_register_file_0_n_38_16), .A1(
      execution_unit_0_register_file_0_n_38_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[15]), .B1(
      execution_unit_0_register_file_0_r6_wr), .B2(pc_sw[15]));
  INV_X1_LVT execution_unit_0_register_file_0_i_38_32 (.ZN(
      execution_unit_0_register_file_0_n_81), .A(
      execution_unit_0_register_file_0_n_38_16));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r6_reg[15] (.Q(
      execution_unit_0_register_file_0_r6[15]), .QN(), .CK(
      execution_unit_0_register_file_0_n_65), .D(
      execution_unit_0_register_file_0_n_81), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_327 (.ZN(
      execution_unit_0_register_file_0_n_105_312), .A1(
      execution_unit_0_register_file_0_n_64), .A2(
      execution_unit_0_register_file_0_r6[15]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_31_31 (.ZN(
      execution_unit_0_register_file_0_n_31_16), .A1(
      execution_unit_0_register_file_0_n_31_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[15]), .B1(
      execution_unit_0_register_file_0_r5_wr), .B2(pc_sw[15]));
  INV_X1_LVT execution_unit_0_register_file_0_i_31_32 (.ZN(
      execution_unit_0_register_file_0_n_62), .A(
      execution_unit_0_register_file_0_n_31_16));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r5_reg[15] (.Q(
      execution_unit_0_register_file_0_r5[15]), .QN(), .CK(
      execution_unit_0_register_file_0_n_46), .D(
      execution_unit_0_register_file_0_n_62), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_328 (.ZN(
      execution_unit_0_register_file_0_n_105_313), .A1(
      execution_unit_0_register_file_0_n_45), .A2(
      execution_unit_0_register_file_0_r5[15]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_105_329 (.ZN(
      execution_unit_0_register_file_0_n_105_314), .A1(
      execution_unit_0_register_file_0_n_105_310), .A2(
      execution_unit_0_register_file_0_n_105_311), .A3(
      execution_unit_0_register_file_0_n_105_312), .A4(
      execution_unit_0_register_file_0_n_105_313));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_87_31 (.ZN(
      execution_unit_0_register_file_0_n_87_16), .A1(
      execution_unit_0_register_file_0_n_87_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[15]), .B1(
      execution_unit_0_register_file_0_r13_wr), .B2(pc_sw[15]));
  INV_X1_LVT execution_unit_0_register_file_0_i_87_32 (.ZN(
      execution_unit_0_register_file_0_n_214), .A(
      execution_unit_0_register_file_0_n_87_16));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r13_reg[15] (.Q(
      execution_unit_0_register_file_0_r13[15]), .QN(), .CK(
      execution_unit_0_register_file_0_n_198), .D(
      execution_unit_0_register_file_0_n_214), .RN(
      execution_unit_0_register_file_0_n_8));
  AND2_X1_LVT execution_unit_0_register_file_0_i_105_330 (.ZN(
      execution_unit_0_register_file_0_n_105_315), .A1(
      execution_unit_0_register_file_0_n_197), .A2(
      execution_unit_0_register_file_0_r13[15]));
  NOR4_X1_LVT execution_unit_0_register_file_0_i_105_331 (.ZN(
      execution_unit_0_register_file_0_n_105_316), .A1(
      execution_unit_0_register_file_0_n_105_304), .A2(
      execution_unit_0_register_file_0_n_105_309), .A3(
      execution_unit_0_register_file_0_n_105_314), .A4(
      execution_unit_0_register_file_0_n_105_315));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_332 (.ZN(
      execution_unit_0_register_file_0_n_105_317), .A1(
      execution_unit_0_register_file_0_n_254), .A2(pc[15]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_101_31 (.ZN(
      execution_unit_0_register_file_0_n_101_16), .A1(
      execution_unit_0_register_file_0_n_101_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[15]), .B1(
      execution_unit_0_register_file_0_r15_wr), .B2(pc_sw[15]));
  INV_X1_LVT execution_unit_0_register_file_0_i_101_32 (.ZN(
      execution_unit_0_register_file_0_n_252), .A(
      execution_unit_0_register_file_0_n_101_16));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r15_reg[15] (.Q(
      execution_unit_0_register_file_0_r15[15]), .QN(), .CK(
      execution_unit_0_register_file_0_n_236), .D(
      execution_unit_0_register_file_0_n_252), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_333 (.ZN(
      execution_unit_0_register_file_0_n_105_318), .A1(
      execution_unit_0_register_file_0_n_235), .A2(
      execution_unit_0_register_file_0_r15[15]));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_94_31 (.ZN(
      execution_unit_0_register_file_0_n_94_16), .A1(
      execution_unit_0_register_file_0_n_94_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[15]), .B1(
      execution_unit_0_register_file_0_r14_wr), .B2(pc_sw[15]));
  INV_X1_LVT execution_unit_0_register_file_0_i_94_32 (.ZN(
      execution_unit_0_register_file_0_n_233), .A(
      execution_unit_0_register_file_0_n_94_16));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r14_reg[15] (.Q(
      execution_unit_0_register_file_0_r14[15]), .QN(), .CK(
      execution_unit_0_register_file_0_n_217), .D(
      execution_unit_0_register_file_0_n_233), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_105_334 (.ZN(
      execution_unit_0_register_file_0_n_105_319), .A1(
      execution_unit_0_register_file_0_n_216), .A2(
      execution_unit_0_register_file_0_r14[15]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_105_335 (.ZN(
      execution_unit_0_reg_src[15]), .A1(
      execution_unit_0_register_file_0_n_105_316), .A2(
      execution_unit_0_register_file_0_n_105_317), .A3(
      execution_unit_0_register_file_0_n_105_318), .A4(
      execution_unit_0_register_file_0_n_105_319));
  XNOR2_X1_LVT execution_unit_0_register_file_0_i_22_15 (.ZN(
      execution_unit_0_register_file_0_n_22_15), .A(execution_unit_0_reg_src[15]), 
      .B(execution_unit_0_register_file_0_n_22_14));
  INV_X1_LVT execution_unit_0_register_file_0_i_22_16 (.ZN(
      execution_unit_0_register_file_0_reg_incr_val[15]), .A(
      execution_unit_0_register_file_0_n_22_15));
  AOI22_X1_LVT execution_unit_0_register_file_0_i_24_31 (.ZN(
      execution_unit_0_register_file_0_n_24_16), .A1(
      execution_unit_0_register_file_0_n_24_0), .A2(
      execution_unit_0_register_file_0_reg_incr_val[15]), .B1(
      execution_unit_0_register_file_0_r4_wr), .B2(pc_sw[15]));
  INV_X1_LVT execution_unit_0_register_file_0_i_24_32 (.ZN(
      execution_unit_0_register_file_0_n_43), .A(
      execution_unit_0_register_file_0_n_24_16));
  DFFR_X1_LVT \execution_unit_0_register_file_0_r4_reg[15] (.Q(
      execution_unit_0_register_file_0_r4[15]), .QN(), .CK(
      execution_unit_0_register_file_0_n_27), .D(
      execution_unit_0_register_file_0_n_43), .RN(
      execution_unit_0_register_file_0_n_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_315 (.ZN(
      execution_unit_0_register_file_0_n_112_300), .A1(inst_dest[4]), .A2(
      execution_unit_0_register_file_0_r4[15]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_316 (.ZN(
      execution_unit_0_register_file_0_n_112_301), .A1(inst_dest[3]), .A2(
      execution_unit_0_register_file_0_r3[15]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_317 (.ZN(
      execution_unit_0_register_file_0_n_112_302), .A1(inst_dest[2]), .A2(
      execution_unit_0_register_file_0_n_0));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_318 (.ZN(
      execution_unit_0_register_file_0_n_112_303), .A1(inst_dest[1]), .A2(
      execution_unit_0_register_file_0_r1[15]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_112_319 (.ZN(
      execution_unit_0_register_file_0_n_112_304), .A1(
      execution_unit_0_register_file_0_n_112_300), .A2(
      execution_unit_0_register_file_0_n_112_301), .A3(
      execution_unit_0_register_file_0_n_112_302), .A4(
      execution_unit_0_register_file_0_n_112_303));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_320 (.ZN(
      execution_unit_0_register_file_0_n_112_305), .A1(inst_dest[12]), .A2(
      execution_unit_0_register_file_0_r12[15]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_321 (.ZN(
      execution_unit_0_register_file_0_n_112_306), .A1(inst_dest[11]), .A2(
      execution_unit_0_register_file_0_r11[15]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_322 (.ZN(
      execution_unit_0_register_file_0_n_112_307), .A1(inst_dest[10]), .A2(
      execution_unit_0_register_file_0_r10[15]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_323 (.ZN(
      execution_unit_0_register_file_0_n_112_308), .A1(inst_dest[9]), .A2(
      execution_unit_0_register_file_0_r9[15]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_112_324 (.ZN(
      execution_unit_0_register_file_0_n_112_309), .A1(
      execution_unit_0_register_file_0_n_112_305), .A2(
      execution_unit_0_register_file_0_n_112_306), .A3(
      execution_unit_0_register_file_0_n_112_307), .A4(
      execution_unit_0_register_file_0_n_112_308));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_325 (.ZN(
      execution_unit_0_register_file_0_n_112_310), .A1(inst_dest[8]), .A2(
      execution_unit_0_register_file_0_r8[15]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_326 (.ZN(
      execution_unit_0_register_file_0_n_112_311), .A1(inst_dest[7]), .A2(
      execution_unit_0_register_file_0_r7[15]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_327 (.ZN(
      execution_unit_0_register_file_0_n_112_312), .A1(inst_dest[6]), .A2(
      execution_unit_0_register_file_0_r6[15]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_328 (.ZN(
      execution_unit_0_register_file_0_n_112_313), .A1(inst_dest[5]), .A2(
      execution_unit_0_register_file_0_r5[15]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_112_329 (.ZN(
      execution_unit_0_register_file_0_n_112_314), .A1(
      execution_unit_0_register_file_0_n_112_310), .A2(
      execution_unit_0_register_file_0_n_112_311), .A3(
      execution_unit_0_register_file_0_n_112_312), .A4(
      execution_unit_0_register_file_0_n_112_313));
  AND2_X1_LVT execution_unit_0_register_file_0_i_112_330 (.ZN(
      execution_unit_0_register_file_0_n_112_315), .A1(inst_dest[13]), .A2(
      execution_unit_0_register_file_0_r13[15]));
  NOR4_X1_LVT execution_unit_0_register_file_0_i_112_331 (.ZN(
      execution_unit_0_register_file_0_n_112_316), .A1(
      execution_unit_0_register_file_0_n_112_304), .A2(
      execution_unit_0_register_file_0_n_112_309), .A3(
      execution_unit_0_register_file_0_n_112_314), .A4(
      execution_unit_0_register_file_0_n_112_315));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_332 (.ZN(
      execution_unit_0_register_file_0_n_112_317), .A1(inst_dest[0]), .A2(pc[15]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_333 (.ZN(
      execution_unit_0_register_file_0_n_112_318), .A1(inst_dest[15]), .A2(
      execution_unit_0_register_file_0_r15[15]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_334 (.ZN(
      execution_unit_0_register_file_0_n_112_319), .A1(inst_dest[14]), .A2(
      execution_unit_0_register_file_0_r14[15]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_112_335 (.ZN(dbg_reg_din[15]), 
      .A1(execution_unit_0_register_file_0_n_112_316), .A2(
      execution_unit_0_register_file_0_n_112_317), .A3(
      execution_unit_0_register_file_0_n_112_318), .A4(
      execution_unit_0_register_file_0_n_112_319));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_294 (.ZN(
      execution_unit_0_register_file_0_n_112_280), .A1(inst_dest[4]), .A2(
      execution_unit_0_register_file_0_r4[14]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_295 (.ZN(
      execution_unit_0_register_file_0_n_112_281), .A1(inst_dest[3]), .A2(
      execution_unit_0_register_file_0_r3[14]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_296 (.ZN(
      execution_unit_0_register_file_0_n_112_282), .A1(inst_dest[2]), .A2(
      execution_unit_0_register_file_0_n_1));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_297 (.ZN(
      execution_unit_0_register_file_0_n_112_283), .A1(inst_dest[1]), .A2(
      execution_unit_0_register_file_0_r1[14]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_112_298 (.ZN(
      execution_unit_0_register_file_0_n_112_284), .A1(
      execution_unit_0_register_file_0_n_112_280), .A2(
      execution_unit_0_register_file_0_n_112_281), .A3(
      execution_unit_0_register_file_0_n_112_282), .A4(
      execution_unit_0_register_file_0_n_112_283));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_299 (.ZN(
      execution_unit_0_register_file_0_n_112_285), .A1(inst_dest[12]), .A2(
      execution_unit_0_register_file_0_r12[14]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_300 (.ZN(
      execution_unit_0_register_file_0_n_112_286), .A1(inst_dest[11]), .A2(
      execution_unit_0_register_file_0_r11[14]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_301 (.ZN(
      execution_unit_0_register_file_0_n_112_287), .A1(inst_dest[10]), .A2(
      execution_unit_0_register_file_0_r10[14]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_302 (.ZN(
      execution_unit_0_register_file_0_n_112_288), .A1(inst_dest[9]), .A2(
      execution_unit_0_register_file_0_r9[14]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_112_303 (.ZN(
      execution_unit_0_register_file_0_n_112_289), .A1(
      execution_unit_0_register_file_0_n_112_285), .A2(
      execution_unit_0_register_file_0_n_112_286), .A3(
      execution_unit_0_register_file_0_n_112_287), .A4(
      execution_unit_0_register_file_0_n_112_288));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_304 (.ZN(
      execution_unit_0_register_file_0_n_112_290), .A1(inst_dest[8]), .A2(
      execution_unit_0_register_file_0_r8[14]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_305 (.ZN(
      execution_unit_0_register_file_0_n_112_291), .A1(inst_dest[7]), .A2(
      execution_unit_0_register_file_0_r7[14]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_306 (.ZN(
      execution_unit_0_register_file_0_n_112_292), .A1(inst_dest[6]), .A2(
      execution_unit_0_register_file_0_r6[14]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_307 (.ZN(
      execution_unit_0_register_file_0_n_112_293), .A1(inst_dest[5]), .A2(
      execution_unit_0_register_file_0_r5[14]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_112_308 (.ZN(
      execution_unit_0_register_file_0_n_112_294), .A1(
      execution_unit_0_register_file_0_n_112_290), .A2(
      execution_unit_0_register_file_0_n_112_291), .A3(
      execution_unit_0_register_file_0_n_112_292), .A4(
      execution_unit_0_register_file_0_n_112_293));
  AND2_X1_LVT execution_unit_0_register_file_0_i_112_309 (.ZN(
      execution_unit_0_register_file_0_n_112_295), .A1(inst_dest[13]), .A2(
      execution_unit_0_register_file_0_r13[14]));
  NOR4_X1_LVT execution_unit_0_register_file_0_i_112_310 (.ZN(
      execution_unit_0_register_file_0_n_112_296), .A1(
      execution_unit_0_register_file_0_n_112_284), .A2(
      execution_unit_0_register_file_0_n_112_289), .A3(
      execution_unit_0_register_file_0_n_112_294), .A4(
      execution_unit_0_register_file_0_n_112_295));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_311 (.ZN(
      execution_unit_0_register_file_0_n_112_297), .A1(inst_dest[0]), .A2(pc[14]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_312 (.ZN(
      execution_unit_0_register_file_0_n_112_298), .A1(inst_dest[15]), .A2(
      execution_unit_0_register_file_0_r15[14]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_313 (.ZN(
      execution_unit_0_register_file_0_n_112_299), .A1(inst_dest[14]), .A2(
      execution_unit_0_register_file_0_r14[14]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_112_314 (.ZN(dbg_reg_din[14]), 
      .A1(execution_unit_0_register_file_0_n_112_296), .A2(
      execution_unit_0_register_file_0_n_112_297), .A3(
      execution_unit_0_register_file_0_n_112_298), .A4(
      execution_unit_0_register_file_0_n_112_299));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_273 (.ZN(
      execution_unit_0_register_file_0_n_112_260), .A1(inst_dest[4]), .A2(
      execution_unit_0_register_file_0_r4[13]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_274 (.ZN(
      execution_unit_0_register_file_0_n_112_261), .A1(inst_dest[3]), .A2(
      execution_unit_0_register_file_0_r3[13]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_275 (.ZN(
      execution_unit_0_register_file_0_n_112_262), .A1(inst_dest[2]), .A2(
      execution_unit_0_register_file_0_n_2));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_276 (.ZN(
      execution_unit_0_register_file_0_n_112_263), .A1(inst_dest[1]), .A2(
      execution_unit_0_register_file_0_r1[13]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_112_277 (.ZN(
      execution_unit_0_register_file_0_n_112_264), .A1(
      execution_unit_0_register_file_0_n_112_260), .A2(
      execution_unit_0_register_file_0_n_112_261), .A3(
      execution_unit_0_register_file_0_n_112_262), .A4(
      execution_unit_0_register_file_0_n_112_263));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_278 (.ZN(
      execution_unit_0_register_file_0_n_112_265), .A1(inst_dest[12]), .A2(
      execution_unit_0_register_file_0_r12[13]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_279 (.ZN(
      execution_unit_0_register_file_0_n_112_266), .A1(inst_dest[11]), .A2(
      execution_unit_0_register_file_0_r11[13]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_280 (.ZN(
      execution_unit_0_register_file_0_n_112_267), .A1(inst_dest[10]), .A2(
      execution_unit_0_register_file_0_r10[13]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_281 (.ZN(
      execution_unit_0_register_file_0_n_112_268), .A1(inst_dest[9]), .A2(
      execution_unit_0_register_file_0_r9[13]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_112_282 (.ZN(
      execution_unit_0_register_file_0_n_112_269), .A1(
      execution_unit_0_register_file_0_n_112_265), .A2(
      execution_unit_0_register_file_0_n_112_266), .A3(
      execution_unit_0_register_file_0_n_112_267), .A4(
      execution_unit_0_register_file_0_n_112_268));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_283 (.ZN(
      execution_unit_0_register_file_0_n_112_270), .A1(inst_dest[8]), .A2(
      execution_unit_0_register_file_0_r8[13]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_284 (.ZN(
      execution_unit_0_register_file_0_n_112_271), .A1(inst_dest[7]), .A2(
      execution_unit_0_register_file_0_r7[13]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_285 (.ZN(
      execution_unit_0_register_file_0_n_112_272), .A1(inst_dest[6]), .A2(
      execution_unit_0_register_file_0_r6[13]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_286 (.ZN(
      execution_unit_0_register_file_0_n_112_273), .A1(inst_dest[5]), .A2(
      execution_unit_0_register_file_0_r5[13]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_112_287 (.ZN(
      execution_unit_0_register_file_0_n_112_274), .A1(
      execution_unit_0_register_file_0_n_112_270), .A2(
      execution_unit_0_register_file_0_n_112_271), .A3(
      execution_unit_0_register_file_0_n_112_272), .A4(
      execution_unit_0_register_file_0_n_112_273));
  AND2_X1_LVT execution_unit_0_register_file_0_i_112_288 (.ZN(
      execution_unit_0_register_file_0_n_112_275), .A1(inst_dest[13]), .A2(
      execution_unit_0_register_file_0_r13[13]));
  NOR4_X1_LVT execution_unit_0_register_file_0_i_112_289 (.ZN(
      execution_unit_0_register_file_0_n_112_276), .A1(
      execution_unit_0_register_file_0_n_112_264), .A2(
      execution_unit_0_register_file_0_n_112_269), .A3(
      execution_unit_0_register_file_0_n_112_274), .A4(
      execution_unit_0_register_file_0_n_112_275));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_290 (.ZN(
      execution_unit_0_register_file_0_n_112_277), .A1(inst_dest[0]), .A2(pc[13]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_291 (.ZN(
      execution_unit_0_register_file_0_n_112_278), .A1(inst_dest[15]), .A2(
      execution_unit_0_register_file_0_r15[13]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_292 (.ZN(
      execution_unit_0_register_file_0_n_112_279), .A1(inst_dest[14]), .A2(
      execution_unit_0_register_file_0_r14[13]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_112_293 (.ZN(dbg_reg_din[13]), 
      .A1(execution_unit_0_register_file_0_n_112_276), .A2(
      execution_unit_0_register_file_0_n_112_277), .A3(
      execution_unit_0_register_file_0_n_112_278), .A4(
      execution_unit_0_register_file_0_n_112_279));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_252 (.ZN(
      execution_unit_0_register_file_0_n_112_240), .A1(inst_dest[4]), .A2(
      execution_unit_0_register_file_0_r4[12]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_253 (.ZN(
      execution_unit_0_register_file_0_n_112_241), .A1(inst_dest[3]), .A2(
      execution_unit_0_register_file_0_r3[12]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_254 (.ZN(
      execution_unit_0_register_file_0_n_112_242), .A1(inst_dest[2]), .A2(
      execution_unit_0_register_file_0_n_3));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_255 (.ZN(
      execution_unit_0_register_file_0_n_112_243), .A1(inst_dest[1]), .A2(
      execution_unit_0_register_file_0_r1[12]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_112_256 (.ZN(
      execution_unit_0_register_file_0_n_112_244), .A1(
      execution_unit_0_register_file_0_n_112_240), .A2(
      execution_unit_0_register_file_0_n_112_241), .A3(
      execution_unit_0_register_file_0_n_112_242), .A4(
      execution_unit_0_register_file_0_n_112_243));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_257 (.ZN(
      execution_unit_0_register_file_0_n_112_245), .A1(inst_dest[12]), .A2(
      execution_unit_0_register_file_0_r12[12]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_258 (.ZN(
      execution_unit_0_register_file_0_n_112_246), .A1(inst_dest[11]), .A2(
      execution_unit_0_register_file_0_r11[12]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_259 (.ZN(
      execution_unit_0_register_file_0_n_112_247), .A1(inst_dest[10]), .A2(
      execution_unit_0_register_file_0_r10[12]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_260 (.ZN(
      execution_unit_0_register_file_0_n_112_248), .A1(inst_dest[9]), .A2(
      execution_unit_0_register_file_0_r9[12]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_112_261 (.ZN(
      execution_unit_0_register_file_0_n_112_249), .A1(
      execution_unit_0_register_file_0_n_112_245), .A2(
      execution_unit_0_register_file_0_n_112_246), .A3(
      execution_unit_0_register_file_0_n_112_247), .A4(
      execution_unit_0_register_file_0_n_112_248));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_262 (.ZN(
      execution_unit_0_register_file_0_n_112_250), .A1(inst_dest[8]), .A2(
      execution_unit_0_register_file_0_r8[12]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_263 (.ZN(
      execution_unit_0_register_file_0_n_112_251), .A1(inst_dest[7]), .A2(
      execution_unit_0_register_file_0_r7[12]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_264 (.ZN(
      execution_unit_0_register_file_0_n_112_252), .A1(inst_dest[6]), .A2(
      execution_unit_0_register_file_0_r6[12]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_265 (.ZN(
      execution_unit_0_register_file_0_n_112_253), .A1(inst_dest[5]), .A2(
      execution_unit_0_register_file_0_r5[12]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_112_266 (.ZN(
      execution_unit_0_register_file_0_n_112_254), .A1(
      execution_unit_0_register_file_0_n_112_250), .A2(
      execution_unit_0_register_file_0_n_112_251), .A3(
      execution_unit_0_register_file_0_n_112_252), .A4(
      execution_unit_0_register_file_0_n_112_253));
  AND2_X1_LVT execution_unit_0_register_file_0_i_112_267 (.ZN(
      execution_unit_0_register_file_0_n_112_255), .A1(inst_dest[13]), .A2(
      execution_unit_0_register_file_0_r13[12]));
  NOR4_X1_LVT execution_unit_0_register_file_0_i_112_268 (.ZN(
      execution_unit_0_register_file_0_n_112_256), .A1(
      execution_unit_0_register_file_0_n_112_244), .A2(
      execution_unit_0_register_file_0_n_112_249), .A3(
      execution_unit_0_register_file_0_n_112_254), .A4(
      execution_unit_0_register_file_0_n_112_255));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_269 (.ZN(
      execution_unit_0_register_file_0_n_112_257), .A1(inst_dest[0]), .A2(pc[12]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_270 (.ZN(
      execution_unit_0_register_file_0_n_112_258), .A1(inst_dest[15]), .A2(
      execution_unit_0_register_file_0_r15[12]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_271 (.ZN(
      execution_unit_0_register_file_0_n_112_259), .A1(inst_dest[14]), .A2(
      execution_unit_0_register_file_0_r14[12]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_112_272 (.ZN(dbg_reg_din[12]), 
      .A1(execution_unit_0_register_file_0_n_112_256), .A2(
      execution_unit_0_register_file_0_n_112_257), .A3(
      execution_unit_0_register_file_0_n_112_258), .A4(
      execution_unit_0_register_file_0_n_112_259));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_231 (.ZN(
      execution_unit_0_register_file_0_n_112_220), .A1(inst_dest[4]), .A2(
      execution_unit_0_register_file_0_r4[11]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_232 (.ZN(
      execution_unit_0_register_file_0_n_112_221), .A1(inst_dest[3]), .A2(
      execution_unit_0_register_file_0_r3[11]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_233 (.ZN(
      execution_unit_0_register_file_0_n_112_222), .A1(inst_dest[2]), .A2(
      execution_unit_0_register_file_0_n_4));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_234 (.ZN(
      execution_unit_0_register_file_0_n_112_223), .A1(inst_dest[1]), .A2(
      execution_unit_0_register_file_0_r1[11]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_112_235 (.ZN(
      execution_unit_0_register_file_0_n_112_224), .A1(
      execution_unit_0_register_file_0_n_112_220), .A2(
      execution_unit_0_register_file_0_n_112_221), .A3(
      execution_unit_0_register_file_0_n_112_222), .A4(
      execution_unit_0_register_file_0_n_112_223));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_236 (.ZN(
      execution_unit_0_register_file_0_n_112_225), .A1(inst_dest[12]), .A2(
      execution_unit_0_register_file_0_r12[11]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_237 (.ZN(
      execution_unit_0_register_file_0_n_112_226), .A1(inst_dest[11]), .A2(
      execution_unit_0_register_file_0_r11[11]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_238 (.ZN(
      execution_unit_0_register_file_0_n_112_227), .A1(inst_dest[10]), .A2(
      execution_unit_0_register_file_0_r10[11]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_239 (.ZN(
      execution_unit_0_register_file_0_n_112_228), .A1(inst_dest[9]), .A2(
      execution_unit_0_register_file_0_r9[11]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_112_240 (.ZN(
      execution_unit_0_register_file_0_n_112_229), .A1(
      execution_unit_0_register_file_0_n_112_225), .A2(
      execution_unit_0_register_file_0_n_112_226), .A3(
      execution_unit_0_register_file_0_n_112_227), .A4(
      execution_unit_0_register_file_0_n_112_228));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_241 (.ZN(
      execution_unit_0_register_file_0_n_112_230), .A1(inst_dest[8]), .A2(
      execution_unit_0_register_file_0_r8[11]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_242 (.ZN(
      execution_unit_0_register_file_0_n_112_231), .A1(inst_dest[7]), .A2(
      execution_unit_0_register_file_0_r7[11]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_243 (.ZN(
      execution_unit_0_register_file_0_n_112_232), .A1(inst_dest[6]), .A2(
      execution_unit_0_register_file_0_r6[11]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_244 (.ZN(
      execution_unit_0_register_file_0_n_112_233), .A1(inst_dest[5]), .A2(
      execution_unit_0_register_file_0_r5[11]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_112_245 (.ZN(
      execution_unit_0_register_file_0_n_112_234), .A1(
      execution_unit_0_register_file_0_n_112_230), .A2(
      execution_unit_0_register_file_0_n_112_231), .A3(
      execution_unit_0_register_file_0_n_112_232), .A4(
      execution_unit_0_register_file_0_n_112_233));
  AND2_X1_LVT execution_unit_0_register_file_0_i_112_246 (.ZN(
      execution_unit_0_register_file_0_n_112_235), .A1(inst_dest[13]), .A2(
      execution_unit_0_register_file_0_r13[11]));
  NOR4_X1_LVT execution_unit_0_register_file_0_i_112_247 (.ZN(
      execution_unit_0_register_file_0_n_112_236), .A1(
      execution_unit_0_register_file_0_n_112_224), .A2(
      execution_unit_0_register_file_0_n_112_229), .A3(
      execution_unit_0_register_file_0_n_112_234), .A4(
      execution_unit_0_register_file_0_n_112_235));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_248 (.ZN(
      execution_unit_0_register_file_0_n_112_237), .A1(inst_dest[0]), .A2(pc[11]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_249 (.ZN(
      execution_unit_0_register_file_0_n_112_238), .A1(inst_dest[15]), .A2(
      execution_unit_0_register_file_0_r15[11]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_250 (.ZN(
      execution_unit_0_register_file_0_n_112_239), .A1(inst_dest[14]), .A2(
      execution_unit_0_register_file_0_r14[11]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_112_251 (.ZN(dbg_reg_din[11]), 
      .A1(execution_unit_0_register_file_0_n_112_236), .A2(
      execution_unit_0_register_file_0_n_112_237), .A3(
      execution_unit_0_register_file_0_n_112_238), .A4(
      execution_unit_0_register_file_0_n_112_239));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_210 (.ZN(
      execution_unit_0_register_file_0_n_112_200), .A1(inst_dest[4]), .A2(
      execution_unit_0_register_file_0_r4[10]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_211 (.ZN(
      execution_unit_0_register_file_0_n_112_201), .A1(inst_dest[3]), .A2(
      execution_unit_0_register_file_0_r3[10]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_212 (.ZN(
      execution_unit_0_register_file_0_n_112_202), .A1(inst_dest[2]), .A2(
      execution_unit_0_register_file_0_n_5));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_213 (.ZN(
      execution_unit_0_register_file_0_n_112_203), .A1(inst_dest[1]), .A2(
      execution_unit_0_register_file_0_r1[10]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_112_214 (.ZN(
      execution_unit_0_register_file_0_n_112_204), .A1(
      execution_unit_0_register_file_0_n_112_200), .A2(
      execution_unit_0_register_file_0_n_112_201), .A3(
      execution_unit_0_register_file_0_n_112_202), .A4(
      execution_unit_0_register_file_0_n_112_203));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_215 (.ZN(
      execution_unit_0_register_file_0_n_112_205), .A1(inst_dest[12]), .A2(
      execution_unit_0_register_file_0_r12[10]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_216 (.ZN(
      execution_unit_0_register_file_0_n_112_206), .A1(inst_dest[11]), .A2(
      execution_unit_0_register_file_0_r11[10]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_217 (.ZN(
      execution_unit_0_register_file_0_n_112_207), .A1(inst_dest[10]), .A2(
      execution_unit_0_register_file_0_r10[10]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_218 (.ZN(
      execution_unit_0_register_file_0_n_112_208), .A1(inst_dest[9]), .A2(
      execution_unit_0_register_file_0_r9[10]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_112_219 (.ZN(
      execution_unit_0_register_file_0_n_112_209), .A1(
      execution_unit_0_register_file_0_n_112_205), .A2(
      execution_unit_0_register_file_0_n_112_206), .A3(
      execution_unit_0_register_file_0_n_112_207), .A4(
      execution_unit_0_register_file_0_n_112_208));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_220 (.ZN(
      execution_unit_0_register_file_0_n_112_210), .A1(inst_dest[8]), .A2(
      execution_unit_0_register_file_0_r8[10]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_221 (.ZN(
      execution_unit_0_register_file_0_n_112_211), .A1(inst_dest[7]), .A2(
      execution_unit_0_register_file_0_r7[10]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_222 (.ZN(
      execution_unit_0_register_file_0_n_112_212), .A1(inst_dest[6]), .A2(
      execution_unit_0_register_file_0_r6[10]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_223 (.ZN(
      execution_unit_0_register_file_0_n_112_213), .A1(inst_dest[5]), .A2(
      execution_unit_0_register_file_0_r5[10]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_112_224 (.ZN(
      execution_unit_0_register_file_0_n_112_214), .A1(
      execution_unit_0_register_file_0_n_112_210), .A2(
      execution_unit_0_register_file_0_n_112_211), .A3(
      execution_unit_0_register_file_0_n_112_212), .A4(
      execution_unit_0_register_file_0_n_112_213));
  AND2_X1_LVT execution_unit_0_register_file_0_i_112_225 (.ZN(
      execution_unit_0_register_file_0_n_112_215), .A1(inst_dest[13]), .A2(
      execution_unit_0_register_file_0_r13[10]));
  NOR4_X1_LVT execution_unit_0_register_file_0_i_112_226 (.ZN(
      execution_unit_0_register_file_0_n_112_216), .A1(
      execution_unit_0_register_file_0_n_112_204), .A2(
      execution_unit_0_register_file_0_n_112_209), .A3(
      execution_unit_0_register_file_0_n_112_214), .A4(
      execution_unit_0_register_file_0_n_112_215));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_227 (.ZN(
      execution_unit_0_register_file_0_n_112_217), .A1(inst_dest[0]), .A2(pc[10]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_228 (.ZN(
      execution_unit_0_register_file_0_n_112_218), .A1(inst_dest[15]), .A2(
      execution_unit_0_register_file_0_r15[10]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_229 (.ZN(
      execution_unit_0_register_file_0_n_112_219), .A1(inst_dest[14]), .A2(
      execution_unit_0_register_file_0_r14[10]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_112_230 (.ZN(dbg_reg_din[10]), 
      .A1(execution_unit_0_register_file_0_n_112_216), .A2(
      execution_unit_0_register_file_0_n_112_217), .A3(
      execution_unit_0_register_file_0_n_112_218), .A4(
      execution_unit_0_register_file_0_n_112_219));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_189 (.ZN(
      execution_unit_0_register_file_0_n_112_180), .A1(inst_dest[4]), .A2(
      execution_unit_0_register_file_0_r4[9]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_190 (.ZN(
      execution_unit_0_register_file_0_n_112_181), .A1(inst_dest[3]), .A2(
      execution_unit_0_register_file_0_r3[9]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_191 (.ZN(
      execution_unit_0_register_file_0_n_112_182), .A1(inst_dest[2]), .A2(
      execution_unit_0_register_file_0_n_6));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_192 (.ZN(
      execution_unit_0_register_file_0_n_112_183), .A1(inst_dest[1]), .A2(
      execution_unit_0_register_file_0_r1[9]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_112_193 (.ZN(
      execution_unit_0_register_file_0_n_112_184), .A1(
      execution_unit_0_register_file_0_n_112_180), .A2(
      execution_unit_0_register_file_0_n_112_181), .A3(
      execution_unit_0_register_file_0_n_112_182), .A4(
      execution_unit_0_register_file_0_n_112_183));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_194 (.ZN(
      execution_unit_0_register_file_0_n_112_185), .A1(inst_dest[12]), .A2(
      execution_unit_0_register_file_0_r12[9]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_195 (.ZN(
      execution_unit_0_register_file_0_n_112_186), .A1(inst_dest[11]), .A2(
      execution_unit_0_register_file_0_r11[9]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_196 (.ZN(
      execution_unit_0_register_file_0_n_112_187), .A1(inst_dest[10]), .A2(
      execution_unit_0_register_file_0_r10[9]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_197 (.ZN(
      execution_unit_0_register_file_0_n_112_188), .A1(inst_dest[9]), .A2(
      execution_unit_0_register_file_0_r9[9]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_112_198 (.ZN(
      execution_unit_0_register_file_0_n_112_189), .A1(
      execution_unit_0_register_file_0_n_112_185), .A2(
      execution_unit_0_register_file_0_n_112_186), .A3(
      execution_unit_0_register_file_0_n_112_187), .A4(
      execution_unit_0_register_file_0_n_112_188));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_199 (.ZN(
      execution_unit_0_register_file_0_n_112_190), .A1(inst_dest[8]), .A2(
      execution_unit_0_register_file_0_r8[9]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_200 (.ZN(
      execution_unit_0_register_file_0_n_112_191), .A1(inst_dest[7]), .A2(
      execution_unit_0_register_file_0_r7[9]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_201 (.ZN(
      execution_unit_0_register_file_0_n_112_192), .A1(inst_dest[6]), .A2(
      execution_unit_0_register_file_0_r6[9]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_202 (.ZN(
      execution_unit_0_register_file_0_n_112_193), .A1(inst_dest[5]), .A2(
      execution_unit_0_register_file_0_r5[9]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_112_203 (.ZN(
      execution_unit_0_register_file_0_n_112_194), .A1(
      execution_unit_0_register_file_0_n_112_190), .A2(
      execution_unit_0_register_file_0_n_112_191), .A3(
      execution_unit_0_register_file_0_n_112_192), .A4(
      execution_unit_0_register_file_0_n_112_193));
  AND2_X1_LVT execution_unit_0_register_file_0_i_112_204 (.ZN(
      execution_unit_0_register_file_0_n_112_195), .A1(inst_dest[13]), .A2(
      execution_unit_0_register_file_0_r13[9]));
  NOR4_X1_LVT execution_unit_0_register_file_0_i_112_205 (.ZN(
      execution_unit_0_register_file_0_n_112_196), .A1(
      execution_unit_0_register_file_0_n_112_184), .A2(
      execution_unit_0_register_file_0_n_112_189), .A3(
      execution_unit_0_register_file_0_n_112_194), .A4(
      execution_unit_0_register_file_0_n_112_195));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_206 (.ZN(
      execution_unit_0_register_file_0_n_112_197), .A1(inst_dest[0]), .A2(pc[9]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_207 (.ZN(
      execution_unit_0_register_file_0_n_112_198), .A1(inst_dest[15]), .A2(
      execution_unit_0_register_file_0_r15[9]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_208 (.ZN(
      execution_unit_0_register_file_0_n_112_199), .A1(inst_dest[14]), .A2(
      execution_unit_0_register_file_0_r14[9]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_112_209 (.ZN(dbg_reg_din[9]), 
      .A1(execution_unit_0_register_file_0_n_112_196), .A2(
      execution_unit_0_register_file_0_n_112_197), .A3(
      execution_unit_0_register_file_0_n_112_198), .A4(
      execution_unit_0_register_file_0_n_112_199));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_168 (.ZN(
      execution_unit_0_register_file_0_n_112_160), .A1(inst_dest[4]), .A2(
      execution_unit_0_register_file_0_r4[8]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_169 (.ZN(
      execution_unit_0_register_file_0_n_112_161), .A1(inst_dest[3]), .A2(
      execution_unit_0_register_file_0_r3[8]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_170 (.ZN(
      execution_unit_0_register_file_0_n_112_162), .A1(inst_dest[2]), .A2(
      execution_unit_0_status[3]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_171 (.ZN(
      execution_unit_0_register_file_0_n_112_163), .A1(inst_dest[1]), .A2(
      execution_unit_0_register_file_0_r1[8]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_112_172 (.ZN(
      execution_unit_0_register_file_0_n_112_164), .A1(
      execution_unit_0_register_file_0_n_112_160), .A2(
      execution_unit_0_register_file_0_n_112_161), .A3(
      execution_unit_0_register_file_0_n_112_162), .A4(
      execution_unit_0_register_file_0_n_112_163));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_173 (.ZN(
      execution_unit_0_register_file_0_n_112_165), .A1(inst_dest[12]), .A2(
      execution_unit_0_register_file_0_r12[8]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_174 (.ZN(
      execution_unit_0_register_file_0_n_112_166), .A1(inst_dest[11]), .A2(
      execution_unit_0_register_file_0_r11[8]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_175 (.ZN(
      execution_unit_0_register_file_0_n_112_167), .A1(inst_dest[10]), .A2(
      execution_unit_0_register_file_0_r10[8]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_176 (.ZN(
      execution_unit_0_register_file_0_n_112_168), .A1(inst_dest[9]), .A2(
      execution_unit_0_register_file_0_r9[8]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_112_177 (.ZN(
      execution_unit_0_register_file_0_n_112_169), .A1(
      execution_unit_0_register_file_0_n_112_165), .A2(
      execution_unit_0_register_file_0_n_112_166), .A3(
      execution_unit_0_register_file_0_n_112_167), .A4(
      execution_unit_0_register_file_0_n_112_168));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_178 (.ZN(
      execution_unit_0_register_file_0_n_112_170), .A1(inst_dest[8]), .A2(
      execution_unit_0_register_file_0_r8[8]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_179 (.ZN(
      execution_unit_0_register_file_0_n_112_171), .A1(inst_dest[7]), .A2(
      execution_unit_0_register_file_0_r7[8]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_180 (.ZN(
      execution_unit_0_register_file_0_n_112_172), .A1(inst_dest[6]), .A2(
      execution_unit_0_register_file_0_r6[8]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_181 (.ZN(
      execution_unit_0_register_file_0_n_112_173), .A1(inst_dest[5]), .A2(
      execution_unit_0_register_file_0_r5[8]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_112_182 (.ZN(
      execution_unit_0_register_file_0_n_112_174), .A1(
      execution_unit_0_register_file_0_n_112_170), .A2(
      execution_unit_0_register_file_0_n_112_171), .A3(
      execution_unit_0_register_file_0_n_112_172), .A4(
      execution_unit_0_register_file_0_n_112_173));
  AND2_X1_LVT execution_unit_0_register_file_0_i_112_183 (.ZN(
      execution_unit_0_register_file_0_n_112_175), .A1(inst_dest[13]), .A2(
      execution_unit_0_register_file_0_r13[8]));
  NOR4_X1_LVT execution_unit_0_register_file_0_i_112_184 (.ZN(
      execution_unit_0_register_file_0_n_112_176), .A1(
      execution_unit_0_register_file_0_n_112_164), .A2(
      execution_unit_0_register_file_0_n_112_169), .A3(
      execution_unit_0_register_file_0_n_112_174), .A4(
      execution_unit_0_register_file_0_n_112_175));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_185 (.ZN(
      execution_unit_0_register_file_0_n_112_177), .A1(inst_dest[0]), .A2(pc[8]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_186 (.ZN(
      execution_unit_0_register_file_0_n_112_178), .A1(inst_dest[15]), .A2(
      execution_unit_0_register_file_0_r15[8]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_187 (.ZN(
      execution_unit_0_register_file_0_n_112_179), .A1(inst_dest[14]), .A2(
      execution_unit_0_register_file_0_r14[8]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_112_188 (.ZN(dbg_reg_din[8]), 
      .A1(execution_unit_0_register_file_0_n_112_176), .A2(
      execution_unit_0_register_file_0_n_112_177), .A3(
      execution_unit_0_register_file_0_n_112_178), .A4(
      execution_unit_0_register_file_0_n_112_179));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_147 (.ZN(
      execution_unit_0_register_file_0_n_112_140), .A1(inst_dest[4]), .A2(
      execution_unit_0_register_file_0_r4[7]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_148 (.ZN(
      execution_unit_0_register_file_0_n_112_141), .A1(inst_dest[3]), .A2(
      execution_unit_0_register_file_0_r3[7]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_149 (.ZN(
      execution_unit_0_register_file_0_n_112_142), .A1(inst_dest[2]), .A2(scg1));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_150 (.ZN(
      execution_unit_0_register_file_0_n_112_143), .A1(inst_dest[1]), .A2(
      execution_unit_0_register_file_0_r1[7]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_112_151 (.ZN(
      execution_unit_0_register_file_0_n_112_144), .A1(
      execution_unit_0_register_file_0_n_112_140), .A2(
      execution_unit_0_register_file_0_n_112_141), .A3(
      execution_unit_0_register_file_0_n_112_142), .A4(
      execution_unit_0_register_file_0_n_112_143));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_152 (.ZN(
      execution_unit_0_register_file_0_n_112_145), .A1(inst_dest[12]), .A2(
      execution_unit_0_register_file_0_r12[7]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_153 (.ZN(
      execution_unit_0_register_file_0_n_112_146), .A1(inst_dest[11]), .A2(
      execution_unit_0_register_file_0_r11[7]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_154 (.ZN(
      execution_unit_0_register_file_0_n_112_147), .A1(inst_dest[10]), .A2(
      execution_unit_0_register_file_0_r10[7]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_155 (.ZN(
      execution_unit_0_register_file_0_n_112_148), .A1(inst_dest[9]), .A2(
      execution_unit_0_register_file_0_r9[7]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_112_156 (.ZN(
      execution_unit_0_register_file_0_n_112_149), .A1(
      execution_unit_0_register_file_0_n_112_145), .A2(
      execution_unit_0_register_file_0_n_112_146), .A3(
      execution_unit_0_register_file_0_n_112_147), .A4(
      execution_unit_0_register_file_0_n_112_148));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_157 (.ZN(
      execution_unit_0_register_file_0_n_112_150), .A1(inst_dest[8]), .A2(
      execution_unit_0_register_file_0_r8[7]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_158 (.ZN(
      execution_unit_0_register_file_0_n_112_151), .A1(inst_dest[7]), .A2(
      execution_unit_0_register_file_0_r7[7]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_159 (.ZN(
      execution_unit_0_register_file_0_n_112_152), .A1(inst_dest[6]), .A2(
      execution_unit_0_register_file_0_r6[7]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_160 (.ZN(
      execution_unit_0_register_file_0_n_112_153), .A1(inst_dest[5]), .A2(
      execution_unit_0_register_file_0_r5[7]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_112_161 (.ZN(
      execution_unit_0_register_file_0_n_112_154), .A1(
      execution_unit_0_register_file_0_n_112_150), .A2(
      execution_unit_0_register_file_0_n_112_151), .A3(
      execution_unit_0_register_file_0_n_112_152), .A4(
      execution_unit_0_register_file_0_n_112_153));
  AND2_X1_LVT execution_unit_0_register_file_0_i_112_162 (.ZN(
      execution_unit_0_register_file_0_n_112_155), .A1(inst_dest[13]), .A2(
      execution_unit_0_register_file_0_r13[7]));
  NOR4_X1_LVT execution_unit_0_register_file_0_i_112_163 (.ZN(
      execution_unit_0_register_file_0_n_112_156), .A1(
      execution_unit_0_register_file_0_n_112_144), .A2(
      execution_unit_0_register_file_0_n_112_149), .A3(
      execution_unit_0_register_file_0_n_112_154), .A4(
      execution_unit_0_register_file_0_n_112_155));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_164 (.ZN(
      execution_unit_0_register_file_0_n_112_157), .A1(inst_dest[0]), .A2(pc[7]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_165 (.ZN(
      execution_unit_0_register_file_0_n_112_158), .A1(inst_dest[15]), .A2(
      execution_unit_0_register_file_0_r15[7]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_166 (.ZN(
      execution_unit_0_register_file_0_n_112_159), .A1(inst_dest[14]), .A2(
      execution_unit_0_register_file_0_r14[7]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_112_167 (.ZN(dbg_reg_din[7]), 
      .A1(execution_unit_0_register_file_0_n_112_156), .A2(
      execution_unit_0_register_file_0_n_112_157), .A3(
      execution_unit_0_register_file_0_n_112_158), .A4(
      execution_unit_0_register_file_0_n_112_159));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_126 (.ZN(
      execution_unit_0_register_file_0_n_112_120), .A1(inst_dest[4]), .A2(
      execution_unit_0_register_file_0_r4[6]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_127 (.ZN(
      execution_unit_0_register_file_0_n_112_121), .A1(inst_dest[3]), .A2(
      execution_unit_0_register_file_0_r3[6]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_128 (.ZN(
      execution_unit_0_register_file_0_n_112_122), .A1(inst_dest[2]), .A2(scg0));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_129 (.ZN(
      execution_unit_0_register_file_0_n_112_123), .A1(inst_dest[1]), .A2(
      execution_unit_0_register_file_0_r1[6]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_112_130 (.ZN(
      execution_unit_0_register_file_0_n_112_124), .A1(
      execution_unit_0_register_file_0_n_112_120), .A2(
      execution_unit_0_register_file_0_n_112_121), .A3(
      execution_unit_0_register_file_0_n_112_122), .A4(
      execution_unit_0_register_file_0_n_112_123));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_131 (.ZN(
      execution_unit_0_register_file_0_n_112_125), .A1(inst_dest[12]), .A2(
      execution_unit_0_register_file_0_r12[6]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_132 (.ZN(
      execution_unit_0_register_file_0_n_112_126), .A1(inst_dest[11]), .A2(
      execution_unit_0_register_file_0_r11[6]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_133 (.ZN(
      execution_unit_0_register_file_0_n_112_127), .A1(inst_dest[10]), .A2(
      execution_unit_0_register_file_0_r10[6]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_134 (.ZN(
      execution_unit_0_register_file_0_n_112_128), .A1(inst_dest[9]), .A2(
      execution_unit_0_register_file_0_r9[6]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_112_135 (.ZN(
      execution_unit_0_register_file_0_n_112_129), .A1(
      execution_unit_0_register_file_0_n_112_125), .A2(
      execution_unit_0_register_file_0_n_112_126), .A3(
      execution_unit_0_register_file_0_n_112_127), .A4(
      execution_unit_0_register_file_0_n_112_128));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_136 (.ZN(
      execution_unit_0_register_file_0_n_112_130), .A1(inst_dest[8]), .A2(
      execution_unit_0_register_file_0_r8[6]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_137 (.ZN(
      execution_unit_0_register_file_0_n_112_131), .A1(inst_dest[7]), .A2(
      execution_unit_0_register_file_0_r7[6]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_138 (.ZN(
      execution_unit_0_register_file_0_n_112_132), .A1(inst_dest[6]), .A2(
      execution_unit_0_register_file_0_r6[6]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_139 (.ZN(
      execution_unit_0_register_file_0_n_112_133), .A1(inst_dest[5]), .A2(
      execution_unit_0_register_file_0_r5[6]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_112_140 (.ZN(
      execution_unit_0_register_file_0_n_112_134), .A1(
      execution_unit_0_register_file_0_n_112_130), .A2(
      execution_unit_0_register_file_0_n_112_131), .A3(
      execution_unit_0_register_file_0_n_112_132), .A4(
      execution_unit_0_register_file_0_n_112_133));
  AND2_X1_LVT execution_unit_0_register_file_0_i_112_141 (.ZN(
      execution_unit_0_register_file_0_n_112_135), .A1(inst_dest[13]), .A2(
      execution_unit_0_register_file_0_r13[6]));
  NOR4_X1_LVT execution_unit_0_register_file_0_i_112_142 (.ZN(
      execution_unit_0_register_file_0_n_112_136), .A1(
      execution_unit_0_register_file_0_n_112_124), .A2(
      execution_unit_0_register_file_0_n_112_129), .A3(
      execution_unit_0_register_file_0_n_112_134), .A4(
      execution_unit_0_register_file_0_n_112_135));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_143 (.ZN(
      execution_unit_0_register_file_0_n_112_137), .A1(inst_dest[0]), .A2(pc[6]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_144 (.ZN(
      execution_unit_0_register_file_0_n_112_138), .A1(inst_dest[15]), .A2(
      execution_unit_0_register_file_0_r15[6]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_145 (.ZN(
      execution_unit_0_register_file_0_n_112_139), .A1(inst_dest[14]), .A2(
      execution_unit_0_register_file_0_r14[6]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_112_146 (.ZN(dbg_reg_din[6]), 
      .A1(execution_unit_0_register_file_0_n_112_136), .A2(
      execution_unit_0_register_file_0_n_112_137), .A3(
      execution_unit_0_register_file_0_n_112_138), .A4(
      execution_unit_0_register_file_0_n_112_139));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_105 (.ZN(
      execution_unit_0_register_file_0_n_112_100), .A1(inst_dest[4]), .A2(
      execution_unit_0_register_file_0_r4[5]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_106 (.ZN(
      execution_unit_0_register_file_0_n_112_101), .A1(inst_dest[3]), .A2(
      execution_unit_0_register_file_0_r3[5]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_107 (.ZN(
      execution_unit_0_register_file_0_n_112_102), .A1(inst_dest[2]), .A2(oscoff));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_108 (.ZN(
      execution_unit_0_register_file_0_n_112_103), .A1(inst_dest[1]), .A2(
      execution_unit_0_register_file_0_r1[5]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_112_109 (.ZN(
      execution_unit_0_register_file_0_n_112_104), .A1(
      execution_unit_0_register_file_0_n_112_100), .A2(
      execution_unit_0_register_file_0_n_112_101), .A3(
      execution_unit_0_register_file_0_n_112_102), .A4(
      execution_unit_0_register_file_0_n_112_103));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_110 (.ZN(
      execution_unit_0_register_file_0_n_112_105), .A1(inst_dest[12]), .A2(
      execution_unit_0_register_file_0_r12[5]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_111 (.ZN(
      execution_unit_0_register_file_0_n_112_106), .A1(inst_dest[11]), .A2(
      execution_unit_0_register_file_0_r11[5]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_112 (.ZN(
      execution_unit_0_register_file_0_n_112_107), .A1(inst_dest[10]), .A2(
      execution_unit_0_register_file_0_r10[5]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_113 (.ZN(
      execution_unit_0_register_file_0_n_112_108), .A1(inst_dest[9]), .A2(
      execution_unit_0_register_file_0_r9[5]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_112_114 (.ZN(
      execution_unit_0_register_file_0_n_112_109), .A1(
      execution_unit_0_register_file_0_n_112_105), .A2(
      execution_unit_0_register_file_0_n_112_106), .A3(
      execution_unit_0_register_file_0_n_112_107), .A4(
      execution_unit_0_register_file_0_n_112_108));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_115 (.ZN(
      execution_unit_0_register_file_0_n_112_110), .A1(inst_dest[8]), .A2(
      execution_unit_0_register_file_0_r8[5]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_116 (.ZN(
      execution_unit_0_register_file_0_n_112_111), .A1(inst_dest[7]), .A2(
      execution_unit_0_register_file_0_r7[5]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_117 (.ZN(
      execution_unit_0_register_file_0_n_112_112), .A1(inst_dest[6]), .A2(
      execution_unit_0_register_file_0_r6[5]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_118 (.ZN(
      execution_unit_0_register_file_0_n_112_113), .A1(inst_dest[5]), .A2(
      execution_unit_0_register_file_0_r5[5]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_112_119 (.ZN(
      execution_unit_0_register_file_0_n_112_114), .A1(
      execution_unit_0_register_file_0_n_112_110), .A2(
      execution_unit_0_register_file_0_n_112_111), .A3(
      execution_unit_0_register_file_0_n_112_112), .A4(
      execution_unit_0_register_file_0_n_112_113));
  AND2_X1_LVT execution_unit_0_register_file_0_i_112_120 (.ZN(
      execution_unit_0_register_file_0_n_112_115), .A1(inst_dest[13]), .A2(
      execution_unit_0_register_file_0_r13[5]));
  NOR4_X1_LVT execution_unit_0_register_file_0_i_112_121 (.ZN(
      execution_unit_0_register_file_0_n_112_116), .A1(
      execution_unit_0_register_file_0_n_112_104), .A2(
      execution_unit_0_register_file_0_n_112_109), .A3(
      execution_unit_0_register_file_0_n_112_114), .A4(
      execution_unit_0_register_file_0_n_112_115));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_122 (.ZN(
      execution_unit_0_register_file_0_n_112_117), .A1(inst_dest[0]), .A2(pc[5]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_123 (.ZN(
      execution_unit_0_register_file_0_n_112_118), .A1(inst_dest[15]), .A2(
      execution_unit_0_register_file_0_r15[5]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_124 (.ZN(
      execution_unit_0_register_file_0_n_112_119), .A1(inst_dest[14]), .A2(
      execution_unit_0_register_file_0_r14[5]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_112_125 (.ZN(dbg_reg_din[5]), 
      .A1(execution_unit_0_register_file_0_n_112_116), .A2(
      execution_unit_0_register_file_0_n_112_117), .A3(
      execution_unit_0_register_file_0_n_112_118), .A4(
      execution_unit_0_register_file_0_n_112_119));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_84 (.ZN(
      execution_unit_0_register_file_0_n_112_80), .A1(inst_dest[4]), .A2(
      execution_unit_0_register_file_0_r4[4]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_85 (.ZN(
      execution_unit_0_register_file_0_n_112_81), .A1(inst_dest[3]), .A2(
      execution_unit_0_register_file_0_r3[4]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_86 (.ZN(
      execution_unit_0_register_file_0_n_112_82), .A1(inst_dest[2]), .A2(
      execution_unit_0_register_file_0_n_7));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_87 (.ZN(
      execution_unit_0_register_file_0_n_112_83), .A1(inst_dest[1]), .A2(
      execution_unit_0_register_file_0_r1[4]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_112_88 (.ZN(
      execution_unit_0_register_file_0_n_112_84), .A1(
      execution_unit_0_register_file_0_n_112_80), .A2(
      execution_unit_0_register_file_0_n_112_81), .A3(
      execution_unit_0_register_file_0_n_112_82), .A4(
      execution_unit_0_register_file_0_n_112_83));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_89 (.ZN(
      execution_unit_0_register_file_0_n_112_85), .A1(inst_dest[12]), .A2(
      execution_unit_0_register_file_0_r12[4]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_90 (.ZN(
      execution_unit_0_register_file_0_n_112_86), .A1(inst_dest[11]), .A2(
      execution_unit_0_register_file_0_r11[4]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_91 (.ZN(
      execution_unit_0_register_file_0_n_112_87), .A1(inst_dest[10]), .A2(
      execution_unit_0_register_file_0_r10[4]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_92 (.ZN(
      execution_unit_0_register_file_0_n_112_88), .A1(inst_dest[9]), .A2(
      execution_unit_0_register_file_0_r9[4]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_112_93 (.ZN(
      execution_unit_0_register_file_0_n_112_89), .A1(
      execution_unit_0_register_file_0_n_112_85), .A2(
      execution_unit_0_register_file_0_n_112_86), .A3(
      execution_unit_0_register_file_0_n_112_87), .A4(
      execution_unit_0_register_file_0_n_112_88));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_94 (.ZN(
      execution_unit_0_register_file_0_n_112_90), .A1(inst_dest[8]), .A2(
      execution_unit_0_register_file_0_r8[4]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_95 (.ZN(
      execution_unit_0_register_file_0_n_112_91), .A1(inst_dest[7]), .A2(
      execution_unit_0_register_file_0_r7[4]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_96 (.ZN(
      execution_unit_0_register_file_0_n_112_92), .A1(inst_dest[6]), .A2(
      execution_unit_0_register_file_0_r6[4]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_97 (.ZN(
      execution_unit_0_register_file_0_n_112_93), .A1(inst_dest[5]), .A2(
      execution_unit_0_register_file_0_r5[4]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_112_98 (.ZN(
      execution_unit_0_register_file_0_n_112_94), .A1(
      execution_unit_0_register_file_0_n_112_90), .A2(
      execution_unit_0_register_file_0_n_112_91), .A3(
      execution_unit_0_register_file_0_n_112_92), .A4(
      execution_unit_0_register_file_0_n_112_93));
  AND2_X1_LVT execution_unit_0_register_file_0_i_112_99 (.ZN(
      execution_unit_0_register_file_0_n_112_95), .A1(inst_dest[13]), .A2(
      execution_unit_0_register_file_0_r13[4]));
  NOR4_X1_LVT execution_unit_0_register_file_0_i_112_100 (.ZN(
      execution_unit_0_register_file_0_n_112_96), .A1(
      execution_unit_0_register_file_0_n_112_84), .A2(
      execution_unit_0_register_file_0_n_112_89), .A3(
      execution_unit_0_register_file_0_n_112_94), .A4(
      execution_unit_0_register_file_0_n_112_95));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_101 (.ZN(
      execution_unit_0_register_file_0_n_112_97), .A1(inst_dest[0]), .A2(pc[4]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_102 (.ZN(
      execution_unit_0_register_file_0_n_112_98), .A1(inst_dest[15]), .A2(
      execution_unit_0_register_file_0_r15[4]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_103 (.ZN(
      execution_unit_0_register_file_0_n_112_99), .A1(inst_dest[14]), .A2(
      execution_unit_0_register_file_0_r14[4]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_112_104 (.ZN(dbg_reg_din[4]), 
      .A1(execution_unit_0_register_file_0_n_112_96), .A2(
      execution_unit_0_register_file_0_n_112_97), .A3(
      execution_unit_0_register_file_0_n_112_98), .A4(
      execution_unit_0_register_file_0_n_112_99));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_63 (.ZN(
      execution_unit_0_register_file_0_n_112_60), .A1(inst_dest[4]), .A2(
      execution_unit_0_register_file_0_r4[3]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_64 (.ZN(
      execution_unit_0_register_file_0_n_112_61), .A1(inst_dest[3]), .A2(
      execution_unit_0_register_file_0_r3[3]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_65 (.ZN(
      execution_unit_0_register_file_0_n_112_62), .A1(inst_dest[2]), .A2(gie));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_66 (.ZN(
      execution_unit_0_register_file_0_n_112_63), .A1(inst_dest[1]), .A2(
      execution_unit_0_register_file_0_r1[3]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_112_67 (.ZN(
      execution_unit_0_register_file_0_n_112_64), .A1(
      execution_unit_0_register_file_0_n_112_60), .A2(
      execution_unit_0_register_file_0_n_112_61), .A3(
      execution_unit_0_register_file_0_n_112_62), .A4(
      execution_unit_0_register_file_0_n_112_63));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_68 (.ZN(
      execution_unit_0_register_file_0_n_112_65), .A1(inst_dest[12]), .A2(
      execution_unit_0_register_file_0_r12[3]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_69 (.ZN(
      execution_unit_0_register_file_0_n_112_66), .A1(inst_dest[11]), .A2(
      execution_unit_0_register_file_0_r11[3]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_70 (.ZN(
      execution_unit_0_register_file_0_n_112_67), .A1(inst_dest[10]), .A2(
      execution_unit_0_register_file_0_r10[3]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_71 (.ZN(
      execution_unit_0_register_file_0_n_112_68), .A1(inst_dest[9]), .A2(
      execution_unit_0_register_file_0_r9[3]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_112_72 (.ZN(
      execution_unit_0_register_file_0_n_112_69), .A1(
      execution_unit_0_register_file_0_n_112_65), .A2(
      execution_unit_0_register_file_0_n_112_66), .A3(
      execution_unit_0_register_file_0_n_112_67), .A4(
      execution_unit_0_register_file_0_n_112_68));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_73 (.ZN(
      execution_unit_0_register_file_0_n_112_70), .A1(inst_dest[8]), .A2(
      execution_unit_0_register_file_0_r8[3]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_74 (.ZN(
      execution_unit_0_register_file_0_n_112_71), .A1(inst_dest[7]), .A2(
      execution_unit_0_register_file_0_r7[3]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_75 (.ZN(
      execution_unit_0_register_file_0_n_112_72), .A1(inst_dest[6]), .A2(
      execution_unit_0_register_file_0_r6[3]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_76 (.ZN(
      execution_unit_0_register_file_0_n_112_73), .A1(inst_dest[5]), .A2(
      execution_unit_0_register_file_0_r5[3]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_112_77 (.ZN(
      execution_unit_0_register_file_0_n_112_74), .A1(
      execution_unit_0_register_file_0_n_112_70), .A2(
      execution_unit_0_register_file_0_n_112_71), .A3(
      execution_unit_0_register_file_0_n_112_72), .A4(
      execution_unit_0_register_file_0_n_112_73));
  AND2_X1_LVT execution_unit_0_register_file_0_i_112_78 (.ZN(
      execution_unit_0_register_file_0_n_112_75), .A1(inst_dest[13]), .A2(
      execution_unit_0_register_file_0_r13[3]));
  NOR4_X1_LVT execution_unit_0_register_file_0_i_112_79 (.ZN(
      execution_unit_0_register_file_0_n_112_76), .A1(
      execution_unit_0_register_file_0_n_112_64), .A2(
      execution_unit_0_register_file_0_n_112_69), .A3(
      execution_unit_0_register_file_0_n_112_74), .A4(
      execution_unit_0_register_file_0_n_112_75));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_80 (.ZN(
      execution_unit_0_register_file_0_n_112_77), .A1(inst_dest[0]), .A2(pc[3]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_81 (.ZN(
      execution_unit_0_register_file_0_n_112_78), .A1(inst_dest[15]), .A2(
      execution_unit_0_register_file_0_r15[3]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_82 (.ZN(
      execution_unit_0_register_file_0_n_112_79), .A1(inst_dest[14]), .A2(
      execution_unit_0_register_file_0_r14[3]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_112_83 (.ZN(dbg_reg_din[3]), 
      .A1(execution_unit_0_register_file_0_n_112_76), .A2(
      execution_unit_0_register_file_0_n_112_77), .A3(
      execution_unit_0_register_file_0_n_112_78), .A4(
      execution_unit_0_register_file_0_n_112_79));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_42 (.ZN(
      execution_unit_0_register_file_0_n_112_40), .A1(inst_dest[4]), .A2(
      execution_unit_0_register_file_0_r4[2]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_43 (.ZN(
      execution_unit_0_register_file_0_n_112_41), .A1(inst_dest[3]), .A2(
      execution_unit_0_register_file_0_r3[2]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_44 (.ZN(
      execution_unit_0_register_file_0_n_112_42), .A1(inst_dest[2]), .A2(
      execution_unit_0_status[2]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_45 (.ZN(
      execution_unit_0_register_file_0_n_112_43), .A1(inst_dest[1]), .A2(
      execution_unit_0_register_file_0_r1[2]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_112_46 (.ZN(
      execution_unit_0_register_file_0_n_112_44), .A1(
      execution_unit_0_register_file_0_n_112_40), .A2(
      execution_unit_0_register_file_0_n_112_41), .A3(
      execution_unit_0_register_file_0_n_112_42), .A4(
      execution_unit_0_register_file_0_n_112_43));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_47 (.ZN(
      execution_unit_0_register_file_0_n_112_45), .A1(inst_dest[12]), .A2(
      execution_unit_0_register_file_0_r12[2]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_48 (.ZN(
      execution_unit_0_register_file_0_n_112_46), .A1(inst_dest[11]), .A2(
      execution_unit_0_register_file_0_r11[2]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_49 (.ZN(
      execution_unit_0_register_file_0_n_112_47), .A1(inst_dest[10]), .A2(
      execution_unit_0_register_file_0_r10[2]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_50 (.ZN(
      execution_unit_0_register_file_0_n_112_48), .A1(inst_dest[9]), .A2(
      execution_unit_0_register_file_0_r9[2]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_112_51 (.ZN(
      execution_unit_0_register_file_0_n_112_49), .A1(
      execution_unit_0_register_file_0_n_112_45), .A2(
      execution_unit_0_register_file_0_n_112_46), .A3(
      execution_unit_0_register_file_0_n_112_47), .A4(
      execution_unit_0_register_file_0_n_112_48));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_52 (.ZN(
      execution_unit_0_register_file_0_n_112_50), .A1(inst_dest[8]), .A2(
      execution_unit_0_register_file_0_r8[2]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_53 (.ZN(
      execution_unit_0_register_file_0_n_112_51), .A1(inst_dest[7]), .A2(
      execution_unit_0_register_file_0_r7[2]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_54 (.ZN(
      execution_unit_0_register_file_0_n_112_52), .A1(inst_dest[6]), .A2(
      execution_unit_0_register_file_0_r6[2]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_55 (.ZN(
      execution_unit_0_register_file_0_n_112_53), .A1(inst_dest[5]), .A2(
      execution_unit_0_register_file_0_r5[2]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_112_56 (.ZN(
      execution_unit_0_register_file_0_n_112_54), .A1(
      execution_unit_0_register_file_0_n_112_50), .A2(
      execution_unit_0_register_file_0_n_112_51), .A3(
      execution_unit_0_register_file_0_n_112_52), .A4(
      execution_unit_0_register_file_0_n_112_53));
  AND2_X1_LVT execution_unit_0_register_file_0_i_112_57 (.ZN(
      execution_unit_0_register_file_0_n_112_55), .A1(inst_dest[13]), .A2(
      execution_unit_0_register_file_0_r13[2]));
  NOR4_X1_LVT execution_unit_0_register_file_0_i_112_58 (.ZN(
      execution_unit_0_register_file_0_n_112_56), .A1(
      execution_unit_0_register_file_0_n_112_44), .A2(
      execution_unit_0_register_file_0_n_112_49), .A3(
      execution_unit_0_register_file_0_n_112_54), .A4(
      execution_unit_0_register_file_0_n_112_55));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_59 (.ZN(
      execution_unit_0_register_file_0_n_112_57), .A1(inst_dest[0]), .A2(pc[2]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_60 (.ZN(
      execution_unit_0_register_file_0_n_112_58), .A1(inst_dest[15]), .A2(
      execution_unit_0_register_file_0_r15[2]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_61 (.ZN(
      execution_unit_0_register_file_0_n_112_59), .A1(inst_dest[14]), .A2(
      execution_unit_0_register_file_0_r14[2]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_112_62 (.ZN(dbg_reg_din[2]), 
      .A1(execution_unit_0_register_file_0_n_112_56), .A2(
      execution_unit_0_register_file_0_n_112_57), .A3(
      execution_unit_0_register_file_0_n_112_58), .A4(
      execution_unit_0_register_file_0_n_112_59));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_21 (.ZN(
      execution_unit_0_register_file_0_n_112_20), .A1(inst_dest[4]), .A2(
      execution_unit_0_register_file_0_r4[1]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_22 (.ZN(
      execution_unit_0_register_file_0_n_112_21), .A1(inst_dest[3]), .A2(
      execution_unit_0_register_file_0_r3[1]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_23 (.ZN(
      execution_unit_0_register_file_0_n_112_22), .A1(inst_dest[2]), .A2(
      execution_unit_0_status[1]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_24 (.ZN(
      execution_unit_0_register_file_0_n_112_23), .A1(inst_dest[1]), .A2(
      execution_unit_0_register_file_0_r1[1]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_112_25 (.ZN(
      execution_unit_0_register_file_0_n_112_24), .A1(
      execution_unit_0_register_file_0_n_112_20), .A2(
      execution_unit_0_register_file_0_n_112_21), .A3(
      execution_unit_0_register_file_0_n_112_22), .A4(
      execution_unit_0_register_file_0_n_112_23));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_26 (.ZN(
      execution_unit_0_register_file_0_n_112_25), .A1(inst_dest[12]), .A2(
      execution_unit_0_register_file_0_r12[1]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_27 (.ZN(
      execution_unit_0_register_file_0_n_112_26), .A1(inst_dest[11]), .A2(
      execution_unit_0_register_file_0_r11[1]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_28 (.ZN(
      execution_unit_0_register_file_0_n_112_27), .A1(inst_dest[10]), .A2(
      execution_unit_0_register_file_0_r10[1]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_29 (.ZN(
      execution_unit_0_register_file_0_n_112_28), .A1(inst_dest[9]), .A2(
      execution_unit_0_register_file_0_r9[1]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_112_30 (.ZN(
      execution_unit_0_register_file_0_n_112_29), .A1(
      execution_unit_0_register_file_0_n_112_25), .A2(
      execution_unit_0_register_file_0_n_112_26), .A3(
      execution_unit_0_register_file_0_n_112_27), .A4(
      execution_unit_0_register_file_0_n_112_28));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_31 (.ZN(
      execution_unit_0_register_file_0_n_112_30), .A1(inst_dest[8]), .A2(
      execution_unit_0_register_file_0_r8[1]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_32 (.ZN(
      execution_unit_0_register_file_0_n_112_31), .A1(inst_dest[7]), .A2(
      execution_unit_0_register_file_0_r7[1]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_33 (.ZN(
      execution_unit_0_register_file_0_n_112_32), .A1(inst_dest[6]), .A2(
      execution_unit_0_register_file_0_r6[1]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_34 (.ZN(
      execution_unit_0_register_file_0_n_112_33), .A1(inst_dest[5]), .A2(
      execution_unit_0_register_file_0_r5[1]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_112_35 (.ZN(
      execution_unit_0_register_file_0_n_112_34), .A1(
      execution_unit_0_register_file_0_n_112_30), .A2(
      execution_unit_0_register_file_0_n_112_31), .A3(
      execution_unit_0_register_file_0_n_112_32), .A4(
      execution_unit_0_register_file_0_n_112_33));
  AND2_X1_LVT execution_unit_0_register_file_0_i_112_36 (.ZN(
      execution_unit_0_register_file_0_n_112_35), .A1(inst_dest[13]), .A2(
      execution_unit_0_register_file_0_r13[1]));
  NOR4_X1_LVT execution_unit_0_register_file_0_i_112_37 (.ZN(
      execution_unit_0_register_file_0_n_112_36), .A1(
      execution_unit_0_register_file_0_n_112_24), .A2(
      execution_unit_0_register_file_0_n_112_29), .A3(
      execution_unit_0_register_file_0_n_112_34), .A4(
      execution_unit_0_register_file_0_n_112_35));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_38 (.ZN(
      execution_unit_0_register_file_0_n_112_37), .A1(inst_dest[0]), .A2(pc[1]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_39 (.ZN(
      execution_unit_0_register_file_0_n_112_38), .A1(inst_dest[15]), .A2(
      execution_unit_0_register_file_0_r15[1]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_40 (.ZN(
      execution_unit_0_register_file_0_n_112_39), .A1(inst_dest[14]), .A2(
      execution_unit_0_register_file_0_r14[1]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_112_41 (.ZN(dbg_reg_din[1]), 
      .A1(execution_unit_0_register_file_0_n_112_36), .A2(
      execution_unit_0_register_file_0_n_112_37), .A3(
      execution_unit_0_register_file_0_n_112_38), .A4(
      execution_unit_0_register_file_0_n_112_39));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_0 (.ZN(
      execution_unit_0_register_file_0_n_112_0), .A1(
      execution_unit_0_register_file_0_r4[0]), .A2(inst_dest[4]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_1 (.ZN(
      execution_unit_0_register_file_0_n_112_1), .A1(
      execution_unit_0_register_file_0_r3[0]), .A2(inst_dest[3]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_2 (.ZN(
      execution_unit_0_register_file_0_n_112_2), .A1(execution_unit_0_status[0]), 
      .A2(inst_dest[2]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_3 (.ZN(
      execution_unit_0_register_file_0_n_112_3), .A1(
      execution_unit_0_register_file_0_r1[0]), .A2(inst_dest[1]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_112_4 (.ZN(
      execution_unit_0_register_file_0_n_112_4), .A1(
      execution_unit_0_register_file_0_n_112_0), .A2(
      execution_unit_0_register_file_0_n_112_1), .A3(
      execution_unit_0_register_file_0_n_112_2), .A4(
      execution_unit_0_register_file_0_n_112_3));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_5 (.ZN(
      execution_unit_0_register_file_0_n_112_5), .A1(
      execution_unit_0_register_file_0_r12[0]), .A2(inst_dest[12]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_6 (.ZN(
      execution_unit_0_register_file_0_n_112_6), .A1(
      execution_unit_0_register_file_0_r11[0]), .A2(inst_dest[11]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_7 (.ZN(
      execution_unit_0_register_file_0_n_112_7), .A1(
      execution_unit_0_register_file_0_r10[0]), .A2(inst_dest[10]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_8 (.ZN(
      execution_unit_0_register_file_0_n_112_8), .A1(
      execution_unit_0_register_file_0_r9[0]), .A2(inst_dest[9]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_112_9 (.ZN(
      execution_unit_0_register_file_0_n_112_9), .A1(
      execution_unit_0_register_file_0_n_112_5), .A2(
      execution_unit_0_register_file_0_n_112_6), .A3(
      execution_unit_0_register_file_0_n_112_7), .A4(
      execution_unit_0_register_file_0_n_112_8));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_10 (.ZN(
      execution_unit_0_register_file_0_n_112_10), .A1(
      execution_unit_0_register_file_0_r8[0]), .A2(inst_dest[8]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_11 (.ZN(
      execution_unit_0_register_file_0_n_112_11), .A1(
      execution_unit_0_register_file_0_r7[0]), .A2(inst_dest[7]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_12 (.ZN(
      execution_unit_0_register_file_0_n_112_12), .A1(
      execution_unit_0_register_file_0_r6[0]), .A2(inst_dest[6]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_13 (.ZN(
      execution_unit_0_register_file_0_n_112_13), .A1(
      execution_unit_0_register_file_0_r5[0]), .A2(inst_dest[5]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_112_14 (.ZN(
      execution_unit_0_register_file_0_n_112_14), .A1(
      execution_unit_0_register_file_0_n_112_10), .A2(
      execution_unit_0_register_file_0_n_112_11), .A3(
      execution_unit_0_register_file_0_n_112_12), .A4(
      execution_unit_0_register_file_0_n_112_13));
  AND2_X1_LVT execution_unit_0_register_file_0_i_112_15 (.ZN(
      execution_unit_0_register_file_0_n_112_15), .A1(
      execution_unit_0_register_file_0_r13[0]), .A2(inst_dest[13]));
  NOR4_X1_LVT execution_unit_0_register_file_0_i_112_16 (.ZN(
      execution_unit_0_register_file_0_n_112_16), .A1(
      execution_unit_0_register_file_0_n_112_4), .A2(
      execution_unit_0_register_file_0_n_112_9), .A3(
      execution_unit_0_register_file_0_n_112_14), .A4(
      execution_unit_0_register_file_0_n_112_15));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_17 (.ZN(
      execution_unit_0_register_file_0_n_112_17), .A1(pc[0]), .A2(inst_dest[0]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_18 (.ZN(
      execution_unit_0_register_file_0_n_112_18), .A1(
      execution_unit_0_register_file_0_r15[0]), .A2(inst_dest[15]));
  NAND2_X1_LVT execution_unit_0_register_file_0_i_112_19 (.ZN(
      execution_unit_0_register_file_0_n_112_19), .A1(
      execution_unit_0_register_file_0_r14[0]), .A2(inst_dest[14]));
  NAND4_X1_LVT execution_unit_0_register_file_0_i_112_20 (.ZN(dbg_reg_din[0]), 
      .A1(execution_unit_0_register_file_0_n_112_16), .A2(
      execution_unit_0_register_file_0_n_112_17), .A3(
      execution_unit_0_register_file_0_n_112_18), .A4(
      execution_unit_0_register_file_0_n_112_19));
  OR2_X1_LVT execution_unit_0_i_8_0 (.ZN(execution_unit_0_n_8_0), .A1(inst_bw), 
      .A2(inst_alu[11]));
  INV_X1_LVT execution_unit_0_i_8_1 (.ZN(execution_unit_0_n_8_1), .A(
      inst_alu[11]));
  NAND2_X1_LVT execution_unit_0_i_8_2 (.ZN(execution_unit_0_n_8_2), .A1(
      execution_unit_0_n_8_1), .A2(inst_bw));
  INV_X1_LVT execution_unit_0_i_8_4 (.ZN(execution_unit_0_n_8_3), .A(eu_mab[0]));
  OAI21_X1_LVT execution_unit_0_i_8_5 (.ZN(execution_unit_0_n_15), .A(
      execution_unit_0_n_8_0), .B1(execution_unit_0_n_8_2), .B2(
      execution_unit_0_n_8_3));
  AND2_X1_LVT execution_unit_0_i_9_1 (.ZN(eu_mb_wr[1]), .A1(
      execution_unit_0_mb_wr_det), .A2(execution_unit_0_n_15));
  OAI21_X1_LVT execution_unit_0_i_8_3 (.ZN(execution_unit_0_n_14), .A(
      execution_unit_0_n_8_0), .B1(execution_unit_0_n_8_2), .B2(eu_mab[0]));
  AND2_X1_LVT execution_unit_0_i_9_0 (.ZN(eu_mb_wr[0]), .A1(
      execution_unit_0_mb_wr_det), .A2(execution_unit_0_n_14));
  INV_X1_LVT execution_unit_0_i_17_0 (.ZN(execution_unit_0_n_17_0), .A(inst_bw));
  NAND2_X1_LVT execution_unit_0_i_13_0 (.ZN(execution_unit_0_n_13_0), .A1(
      e_state[0]), .A2(e_state[3]));
  NOR3_X1_LVT execution_unit_0_i_13_1 (.ZN(execution_unit_0_n_13_1), .A1(
      execution_unit_0_n_13_0), .A2(e_state[1]), .A3(e_state[2]));
  INV_X1_LVT execution_unit_0_i_13_2 (.ZN(execution_unit_0_n_13_2), .A(
      execution_unit_0_n_13_1));
  AOI22_X1_LVT execution_unit_0_i_13_33 (.ZN(execution_unit_0_n_13_18), .A1(
      execution_unit_0_n_13_2), .A2(execution_unit_0_alu_out[15]), .B1(
      execution_unit_0_n_13_1), .B2(pc_nxt[15]));
  INV_X1_LVT execution_unit_0_i_13_34 (.ZN(execution_unit_0_n_34), .A(
      execution_unit_0_n_13_18));
  INV_X1_LVT execution_unit_0_i_14_0 (.ZN(execution_unit_0_n_14_0), .A(
      inst_so[5]));
  AOI211_X1_LVT execution_unit_0_i_14_1 (.ZN(execution_unit_0_n_14_1), .A(
      execution_unit_0_n_7), .B(execution_unit_0_reg_sr_clr), .C1(
      execution_unit_0_n_14_0), .C2(execution_unit_0_n_0));
  INV_X1_LVT execution_unit_0_i_14_2 (.ZN(execution_unit_0_n_35), .A(
      execution_unit_0_n_14_1));
  INV_X1_LVT execution_unit_0_i_15_3 (.ZN(execution_unit_0_n_15_3), .A(
      execution_unit_0_n_35));
  NAND2_X1_LVT execution_unit_0_i_15_0 (.ZN(execution_unit_0_n_15_0), .A1(
      e_state[0]), .A2(e_state[3]));
  NOR3_X1_LVT execution_unit_0_i_15_1 (.ZN(execution_unit_0_n_15_1), .A1(
      execution_unit_0_n_15_0), .A2(e_state[1]), .A3(e_state[2]));
  INV_X1_LVT execution_unit_0_i_15_2 (.ZN(execution_unit_0_n_15_2), .A(
      execution_unit_0_n_15_1));
  NAND2_X1_LVT execution_unit_0_i_15_4 (.ZN(execution_unit_0_n_36), .A1(
      execution_unit_0_n_15_3), .A2(execution_unit_0_n_15_2));
  CLKGATETST_X1_LVT execution_unit_0_clk_gate_mdb_out_nxt_reg (.GCK(
      execution_unit_0_n_17), .CK(cpu_mclk), .E(execution_unit_0_n_36), .SE(1'b0));
  DFFR_X1_LVT \execution_unit_0_mdb_out_nxt_reg[15] (.Q(
      execution_unit_0_mdb_out_nxt[15]), .QN(), .CK(execution_unit_0_n_17), .D(
      execution_unit_0_n_34), .RN(execution_unit_0_n_18));
  AOI22_X1_LVT execution_unit_0_i_13_17 (.ZN(execution_unit_0_n_13_10), .A1(
      execution_unit_0_n_13_2), .A2(execution_unit_0_alu_out[7]), .B1(
      execution_unit_0_n_13_1), .B2(pc_nxt[7]));
  INV_X1_LVT execution_unit_0_i_13_18 (.ZN(execution_unit_0_n_26), .A(
      execution_unit_0_n_13_10));
  DFFR_X1_LVT \execution_unit_0_mdb_out_nxt_reg[7] (.Q(eu_mdb_out[7]), .QN(), 
      .CK(execution_unit_0_n_17), .D(execution_unit_0_n_26), .RN(
      execution_unit_0_n_18));
  AOI22_X1_LVT execution_unit_0_i_17_15 (.ZN(execution_unit_0_n_17_8), .A1(
      execution_unit_0_n_17_0), .A2(execution_unit_0_mdb_out_nxt[15]), .B1(
      inst_bw), .B2(eu_mdb_out[7]));
  INV_X1_LVT execution_unit_0_i_17_16 (.ZN(eu_mdb_out[15]), .A(
      execution_unit_0_n_17_8));
  AOI22_X1_LVT execution_unit_0_i_13_31 (.ZN(execution_unit_0_n_13_17), .A1(
      execution_unit_0_n_13_2), .A2(execution_unit_0_alu_out[14]), .B1(
      execution_unit_0_n_13_1), .B2(pc_nxt[14]));
  INV_X1_LVT execution_unit_0_i_13_32 (.ZN(execution_unit_0_n_33), .A(
      execution_unit_0_n_13_17));
  DFFR_X1_LVT \execution_unit_0_mdb_out_nxt_reg[14] (.Q(
      execution_unit_0_mdb_out_nxt[14]), .QN(), .CK(execution_unit_0_n_17), .D(
      execution_unit_0_n_33), .RN(execution_unit_0_n_18));
  AOI22_X1_LVT execution_unit_0_i_13_15 (.ZN(execution_unit_0_n_13_9), .A1(
      execution_unit_0_n_13_2), .A2(execution_unit_0_alu_out[6]), .B1(
      execution_unit_0_n_13_1), .B2(pc_nxt[6]));
  INV_X1_LVT execution_unit_0_i_13_16 (.ZN(execution_unit_0_n_25), .A(
      execution_unit_0_n_13_9));
  DFFR_X1_LVT \execution_unit_0_mdb_out_nxt_reg[6] (.Q(eu_mdb_out[6]), .QN(), 
      .CK(execution_unit_0_n_17), .D(execution_unit_0_n_25), .RN(
      execution_unit_0_n_18));
  AOI22_X1_LVT execution_unit_0_i_17_13 (.ZN(execution_unit_0_n_17_7), .A1(
      execution_unit_0_n_17_0), .A2(execution_unit_0_mdb_out_nxt[14]), .B1(
      inst_bw), .B2(eu_mdb_out[6]));
  INV_X1_LVT execution_unit_0_i_17_14 (.ZN(eu_mdb_out[14]), .A(
      execution_unit_0_n_17_7));
  AOI22_X1_LVT execution_unit_0_i_13_29 (.ZN(execution_unit_0_n_13_16), .A1(
      execution_unit_0_n_13_2), .A2(execution_unit_0_alu_out[13]), .B1(
      execution_unit_0_n_13_1), .B2(pc_nxt[13]));
  INV_X1_LVT execution_unit_0_i_13_30 (.ZN(execution_unit_0_n_32), .A(
      execution_unit_0_n_13_16));
  DFFR_X1_LVT \execution_unit_0_mdb_out_nxt_reg[13] (.Q(
      execution_unit_0_mdb_out_nxt[13]), .QN(), .CK(execution_unit_0_n_17), .D(
      execution_unit_0_n_32), .RN(execution_unit_0_n_18));
  AOI22_X1_LVT execution_unit_0_i_13_13 (.ZN(execution_unit_0_n_13_8), .A1(
      execution_unit_0_n_13_2), .A2(execution_unit_0_alu_out[5]), .B1(
      execution_unit_0_n_13_1), .B2(pc_nxt[5]));
  INV_X1_LVT execution_unit_0_i_13_14 (.ZN(execution_unit_0_n_24), .A(
      execution_unit_0_n_13_8));
  DFFR_X1_LVT \execution_unit_0_mdb_out_nxt_reg[5] (.Q(eu_mdb_out[5]), .QN(), 
      .CK(execution_unit_0_n_17), .D(execution_unit_0_n_24), .RN(
      execution_unit_0_n_18));
  AOI22_X1_LVT execution_unit_0_i_17_11 (.ZN(execution_unit_0_n_17_6), .A1(
      execution_unit_0_n_17_0), .A2(execution_unit_0_mdb_out_nxt[13]), .B1(
      inst_bw), .B2(eu_mdb_out[5]));
  INV_X1_LVT execution_unit_0_i_17_12 (.ZN(eu_mdb_out[13]), .A(
      execution_unit_0_n_17_6));
  AOI22_X1_LVT execution_unit_0_i_13_27 (.ZN(execution_unit_0_n_13_15), .A1(
      execution_unit_0_n_13_2), .A2(execution_unit_0_alu_out[12]), .B1(
      execution_unit_0_n_13_1), .B2(pc_nxt[12]));
  INV_X1_LVT execution_unit_0_i_13_28 (.ZN(execution_unit_0_n_31), .A(
      execution_unit_0_n_13_15));
  DFFR_X1_LVT \execution_unit_0_mdb_out_nxt_reg[12] (.Q(
      execution_unit_0_mdb_out_nxt[12]), .QN(), .CK(execution_unit_0_n_17), .D(
      execution_unit_0_n_31), .RN(execution_unit_0_n_18));
  AOI22_X1_LVT execution_unit_0_i_13_11 (.ZN(execution_unit_0_n_13_7), .A1(
      execution_unit_0_n_13_2), .A2(execution_unit_0_alu_out[4]), .B1(
      execution_unit_0_n_13_1), .B2(pc_nxt[4]));
  INV_X1_LVT execution_unit_0_i_13_12 (.ZN(execution_unit_0_n_23), .A(
      execution_unit_0_n_13_7));
  DFFR_X1_LVT \execution_unit_0_mdb_out_nxt_reg[4] (.Q(eu_mdb_out[4]), .QN(), 
      .CK(execution_unit_0_n_17), .D(execution_unit_0_n_23), .RN(
      execution_unit_0_n_18));
  AOI22_X1_LVT execution_unit_0_i_17_9 (.ZN(execution_unit_0_n_17_5), .A1(
      execution_unit_0_n_17_0), .A2(execution_unit_0_mdb_out_nxt[12]), .B1(
      inst_bw), .B2(eu_mdb_out[4]));
  INV_X1_LVT execution_unit_0_i_17_10 (.ZN(eu_mdb_out[12]), .A(
      execution_unit_0_n_17_5));
  AOI22_X1_LVT execution_unit_0_i_13_25 (.ZN(execution_unit_0_n_13_14), .A1(
      execution_unit_0_n_13_2), .A2(execution_unit_0_alu_out[11]), .B1(
      execution_unit_0_n_13_1), .B2(pc_nxt[11]));
  INV_X1_LVT execution_unit_0_i_13_26 (.ZN(execution_unit_0_n_30), .A(
      execution_unit_0_n_13_14));
  DFFR_X1_LVT \execution_unit_0_mdb_out_nxt_reg[11] (.Q(
      execution_unit_0_mdb_out_nxt[11]), .QN(), .CK(execution_unit_0_n_17), .D(
      execution_unit_0_n_30), .RN(execution_unit_0_n_18));
  AOI22_X1_LVT execution_unit_0_i_13_9 (.ZN(execution_unit_0_n_13_6), .A1(
      execution_unit_0_n_13_2), .A2(execution_unit_0_alu_out[3]), .B1(
      execution_unit_0_n_13_1), .B2(pc_nxt[3]));
  INV_X1_LVT execution_unit_0_i_13_10 (.ZN(execution_unit_0_n_22), .A(
      execution_unit_0_n_13_6));
  DFFR_X1_LVT \execution_unit_0_mdb_out_nxt_reg[3] (.Q(eu_mdb_out[3]), .QN(), 
      .CK(execution_unit_0_n_17), .D(execution_unit_0_n_22), .RN(
      execution_unit_0_n_18));
  AOI22_X1_LVT execution_unit_0_i_17_7 (.ZN(execution_unit_0_n_17_4), .A1(
      execution_unit_0_n_17_0), .A2(execution_unit_0_mdb_out_nxt[11]), .B1(
      inst_bw), .B2(eu_mdb_out[3]));
  INV_X1_LVT execution_unit_0_i_17_8 (.ZN(eu_mdb_out[11]), .A(
      execution_unit_0_n_17_4));
  AOI22_X1_LVT execution_unit_0_i_13_23 (.ZN(execution_unit_0_n_13_13), .A1(
      execution_unit_0_n_13_2), .A2(execution_unit_0_alu_out[10]), .B1(
      execution_unit_0_n_13_1), .B2(pc_nxt[10]));
  INV_X1_LVT execution_unit_0_i_13_24 (.ZN(execution_unit_0_n_29), .A(
      execution_unit_0_n_13_13));
  DFFR_X1_LVT \execution_unit_0_mdb_out_nxt_reg[10] (.Q(
      execution_unit_0_mdb_out_nxt[10]), .QN(), .CK(execution_unit_0_n_17), .D(
      execution_unit_0_n_29), .RN(execution_unit_0_n_18));
  AOI22_X1_LVT execution_unit_0_i_13_7 (.ZN(execution_unit_0_n_13_5), .A1(
      execution_unit_0_n_13_2), .A2(execution_unit_0_alu_out[2]), .B1(
      execution_unit_0_n_13_1), .B2(pc_nxt[2]));
  INV_X1_LVT execution_unit_0_i_13_8 (.ZN(execution_unit_0_n_21), .A(
      execution_unit_0_n_13_5));
  DFFR_X1_LVT \execution_unit_0_mdb_out_nxt_reg[2] (.Q(eu_mdb_out[2]), .QN(), 
      .CK(execution_unit_0_n_17), .D(execution_unit_0_n_21), .RN(
      execution_unit_0_n_18));
  AOI22_X1_LVT execution_unit_0_i_17_5 (.ZN(execution_unit_0_n_17_3), .A1(
      execution_unit_0_n_17_0), .A2(execution_unit_0_mdb_out_nxt[10]), .B1(
      inst_bw), .B2(eu_mdb_out[2]));
  INV_X1_LVT execution_unit_0_i_17_6 (.ZN(eu_mdb_out[10]), .A(
      execution_unit_0_n_17_3));
  AOI22_X1_LVT execution_unit_0_i_13_21 (.ZN(execution_unit_0_n_13_12), .A1(
      execution_unit_0_n_13_2), .A2(execution_unit_0_alu_out[9]), .B1(
      execution_unit_0_n_13_1), .B2(pc_nxt[9]));
  INV_X1_LVT execution_unit_0_i_13_22 (.ZN(execution_unit_0_n_28), .A(
      execution_unit_0_n_13_12));
  DFFR_X1_LVT \execution_unit_0_mdb_out_nxt_reg[9] (.Q(
      execution_unit_0_mdb_out_nxt[9]), .QN(), .CK(execution_unit_0_n_17), .D(
      execution_unit_0_n_28), .RN(execution_unit_0_n_18));
  AOI22_X1_LVT execution_unit_0_i_13_5 (.ZN(execution_unit_0_n_13_4), .A1(
      execution_unit_0_n_13_2), .A2(execution_unit_0_alu_out[1]), .B1(
      execution_unit_0_n_13_1), .B2(pc_nxt[1]));
  INV_X1_LVT execution_unit_0_i_13_6 (.ZN(execution_unit_0_n_20), .A(
      execution_unit_0_n_13_4));
  DFFR_X1_LVT \execution_unit_0_mdb_out_nxt_reg[1] (.Q(eu_mdb_out[1]), .QN(), 
      .CK(execution_unit_0_n_17), .D(execution_unit_0_n_20), .RN(
      execution_unit_0_n_18));
  AOI22_X1_LVT execution_unit_0_i_17_3 (.ZN(execution_unit_0_n_17_2), .A1(
      execution_unit_0_n_17_0), .A2(execution_unit_0_mdb_out_nxt[9]), .B1(
      inst_bw), .B2(eu_mdb_out[1]));
  INV_X1_LVT execution_unit_0_i_17_4 (.ZN(eu_mdb_out[9]), .A(
      execution_unit_0_n_17_2));
  AOI22_X1_LVT execution_unit_0_i_13_19 (.ZN(execution_unit_0_n_13_11), .A1(
      execution_unit_0_n_13_2), .A2(execution_unit_0_alu_out[8]), .B1(
      execution_unit_0_n_13_1), .B2(pc_nxt[8]));
  INV_X1_LVT execution_unit_0_i_13_20 (.ZN(execution_unit_0_n_27), .A(
      execution_unit_0_n_13_11));
  DFFR_X1_LVT \execution_unit_0_mdb_out_nxt_reg[8] (.Q(
      execution_unit_0_mdb_out_nxt[8]), .QN(), .CK(execution_unit_0_n_17), .D(
      execution_unit_0_n_27), .RN(execution_unit_0_n_18));
  AOI22_X1_LVT execution_unit_0_i_13_3 (.ZN(execution_unit_0_n_13_3), .A1(
      execution_unit_0_n_13_2), .A2(execution_unit_0_alu_out[0]), .B1(
      execution_unit_0_n_13_1), .B2(pc_nxt[0]));
  INV_X1_LVT execution_unit_0_i_13_4 (.ZN(execution_unit_0_n_19), .A(
      execution_unit_0_n_13_3));
  DFFR_X1_LVT \execution_unit_0_mdb_out_nxt_reg[0] (.Q(eu_mdb_out[0]), .QN(), .CK(
      execution_unit_0_n_17), .D(execution_unit_0_n_19), .RN(
      execution_unit_0_n_18));
  AOI22_X1_LVT execution_unit_0_i_17_1 (.ZN(execution_unit_0_n_17_1), .A1(
      execution_unit_0_n_17_0), .A2(execution_unit_0_mdb_out_nxt[8]), .B1(
      eu_mdb_out[0]), .B2(inst_bw));
  INV_X1_LVT execution_unit_0_i_17_2 (.ZN(eu_mdb_out[8]), .A(
      execution_unit_0_n_17_1));
  NAND3_X1_LVT clock_module_0_i_7_0 (.ZN(clock_module_0_n_7_0), .A1(per_addr[3]), 
      .A2(per_addr[5]), .A3(per_en));
  NOR4_X1_LVT clock_module_0_i_7_1 (.ZN(clock_module_0_n_7_1), .A1(
      clock_module_0_n_7_0), .A2(per_addr[11]), .A3(per_addr[12]), .A4(
      per_addr[13]));
  NOR4_X1_LVT clock_module_0_i_7_2 (.ZN(clock_module_0_n_7_2), .A1(per_addr[7]), 
      .A2(per_addr[8]), .A3(per_addr[9]), .A4(per_addr[10]));
  NAND2_X1_LVT clock_module_0_i_7_3 (.ZN(clock_module_0_n_7_3), .A1(
      clock_module_0_n_7_1), .A2(clock_module_0_n_7_2));
  NOR3_X1_LVT clock_module_0_i_7_4 (.ZN(clock_module_0_reg_sel), .A1(
      clock_module_0_n_7_3), .A2(per_addr[4]), .A3(per_addr[6]));
  AND2_X1_LVT clock_module_0_i_16_0 (.ZN(clock_module_0_reg_hi_write), .A1(
      per_we[1]), .A2(clock_module_0_reg_sel));
  NAND2_X1_LVT clock_module_0_i_11_0 (.ZN(clock_module_0_n_11_0), .A1(per_addr[0]), 
      .A2(per_addr[1]));
  NOR2_X1_LVT clock_module_0_i_11_1 (.ZN(clock_module_0_n_5), .A1(
      clock_module_0_n_11_0), .A2(per_addr[2]));
  AND2_X1_LVT clock_module_0_i_17_0 (.ZN(clock_module_0_bcsctl1_wr), .A1(
      clock_module_0_reg_hi_write), .A2(clock_module_0_n_5));
  INV_X1_LVT clock_module_0_i_40_0 (.ZN(clock_module_0_por_a), .A(reset_n));
  INV_X1_LVT clock_module_0_sync_cell_mclk_wkup_i_0_0 (.ZN(
      clock_module_0_sync_cell_mclk_wkup_n_0), .A(puc_rst));
  DFFR_X1_LVT \clock_module_0_sync_cell_mclk_wkup_data_sync_reg[0] (.Q(
      clock_module_0_sync_cell_mclk_wkup_n_1), .QN(), .CK(dco_clk), .D(mclk_wkup), 
      .RN(clock_module_0_sync_cell_mclk_wkup_n_0));
  DFFR_X1_LVT \clock_module_0_sync_cell_mclk_wkup_data_sync_reg[1] (.Q(
      clock_module_0_mclk_wkup_s), .QN(), .CK(dco_clk), .D(
      clock_module_0_sync_cell_mclk_wkup_n_1), .RN(
      clock_module_0_sync_cell_mclk_wkup_n_0));
  NOR2_X1_LVT clock_module_0_i_37_0 (.ZN(clock_module_0_n_37_0), .A1(mclk_enable), 
      .A2(clock_module_0_mclk_wkup_s));
  NAND2_X1_LVT clock_module_0_i_37_1 (.ZN(clock_module_0_n_37_1), .A1(dbg_en), 
      .A2(cpu_en));
  NAND2_X1_LVT clock_module_0_i_37_2 (.ZN(clock_module_0_mclk_active), .A1(
      clock_module_0_n_37_0), .A2(clock_module_0_n_37_1));
  AND2_X1_LVT clock_module_0_i_13_0 (.ZN(clock_module_0_reg_lo_write), .A1(
      per_we[0]), .A2(clock_module_0_reg_sel));
  INV_X1_LVT clock_module_0_i_10_0 (.ZN(clock_module_0_n_10_0), .A(per_addr[2]));
  NOR3_X1_LVT clock_module_0_i_10_1 (.ZN(clock_module_0_n_4), .A1(
      clock_module_0_n_10_0), .A2(per_addr[0]), .A3(per_addr[1]));
  AND2_X1_LVT clock_module_0_i_14_0 (.ZN(clock_module_0_bcsctl2_wr), .A1(
      clock_module_0_reg_lo_write), .A2(clock_module_0_n_4));
  CLKGATETST_X1_LVT clock_module_0_clk_gate_bcsctl2_reg (.GCK(clock_module_0_n_8), 
      .CK(mclk), .E(clock_module_0_bcsctl2_wr), .SE(1'b0));
  DFFR_X1_LVT \clock_module_0_bcsctl2_reg[5] (.Q(clock_module_0_bcsctl2[5]), .QN(), 
      .CK(clock_module_0_n_8), .D(per_din[5]), .RN(clock_module_0_n_10));
  INV_X1_LVT clock_module_0_i_36_2 (.ZN(clock_module_0_n_36_2), .A(
      clock_module_0_bcsctl2[5]));
  DFFR_X1_LVT \clock_module_0_bcsctl2_reg[4] (.Q(clock_module_0_bcsctl2[4]), .QN(), 
      .CK(clock_module_0_n_8), .D(per_din[4]), .RN(clock_module_0_n_10));
  OR2_X1_LVT clock_module_0_i_36_3 (.ZN(clock_module_0_n_36_3), .A1(
      clock_module_0_n_36_2), .A2(clock_module_0_bcsctl2[4]));
  INV_X1_LVT clock_module_0_i_31_0 (.ZN(clock_module_0_n_19), .A(
      clock_module_0_mclk_div[0]));
  OR2_X1_LVT clock_module_0_i_32_0 (.ZN(clock_module_0_n_22), .A1(
      clock_module_0_bcsctl2[4]), .A2(clock_module_0_bcsctl2[5]));
  CLKGATETST_X1_LVT clock_module_0_clk_gate_mclk_div_reg (.GCK(
      clock_module_0_n_18), .CK(dco_clk), .E(clock_module_0_n_22), .SE(1'b0));
  DFFR_X1_LVT \clock_module_0_mclk_div_reg[0] (.Q(clock_module_0_mclk_div[0]), 
      .QN(), .CK(clock_module_0_n_18), .D(clock_module_0_n_19), .RN(
      clock_module_0_n_10));
  HA_X1_LVT clock_module_0_i_31_1 (.CO(clock_module_0_n_31_0), .S(
      clock_module_0_n_20), .A(clock_module_0_mclk_div[1]), .B(
      clock_module_0_mclk_div[0]));
  DFFR_X1_LVT \clock_module_0_mclk_div_reg[1] (.Q(clock_module_0_mclk_div[1]), 
      .QN(), .CK(clock_module_0_n_18), .D(clock_module_0_n_20), .RN(
      clock_module_0_n_10));
  XNOR2_X1_LVT clock_module_0_i_31_2 (.ZN(clock_module_0_n_31_1), .A(
      clock_module_0_mclk_div[2]), .B(clock_module_0_n_31_0));
  INV_X1_LVT clock_module_0_i_31_3 (.ZN(clock_module_0_n_21), .A(
      clock_module_0_n_31_1));
  DFFR_X1_LVT \clock_module_0_mclk_div_reg[2] (.Q(clock_module_0_mclk_div[2]), 
      .QN(), .CK(clock_module_0_n_18), .D(clock_module_0_n_21), .RN(
      clock_module_0_n_10));
  AND3_X1_LVT clock_module_0_i_34_0 (.ZN(clock_module_0_n_23), .A1(
      clock_module_0_mclk_div[0]), .A2(clock_module_0_mclk_div[1]), .A3(
      clock_module_0_mclk_div[2]));
  INV_X1_LVT clock_module_0_i_36_4 (.ZN(clock_module_0_n_36_4), .A(
      clock_module_0_n_36_3));
  AND2_X1_LVT clock_module_0_i_35_0 (.ZN(clock_module_0_n_24), .A1(
      clock_module_0_mclk_div[0]), .A2(clock_module_0_mclk_div[1]));
  AOI22_X1_LVT clock_module_0_i_36_5 (.ZN(clock_module_0_n_36_5), .A1(
      clock_module_0_n_36_3), .A2(clock_module_0_n_23), .B1(
      clock_module_0_n_36_4), .B2(clock_module_0_n_24));
  INV_X1_LVT clock_module_0_i_36_6 (.ZN(clock_module_0_n_36_6), .A(
      clock_module_0_n_36_5));
  NAND2_X1_LVT clock_module_0_i_36_7 (.ZN(clock_module_0_n_36_7), .A1(
      clock_module_0_n_36_2), .A2(clock_module_0_bcsctl2[4]));
  INV_X1_LVT clock_module_0_i_36_8 (.ZN(clock_module_0_n_36_8), .A(
      clock_module_0_n_36_7));
  AOI22_X1_LVT clock_module_0_i_36_9 (.ZN(clock_module_0_n_36_9), .A1(
      clock_module_0_n_36_6), .A2(clock_module_0_n_36_7), .B1(
      clock_module_0_n_36_8), .B2(clock_module_0_mclk_div[0]));
  NOR2_X1_LVT clock_module_0_i_36_0 (.ZN(clock_module_0_n_36_0), .A1(
      clock_module_0_bcsctl2[4]), .A2(clock_module_0_bcsctl2[5]));
  INV_X1_LVT clock_module_0_i_36_1 (.ZN(clock_module_0_n_36_1), .A(
      clock_module_0_n_36_0));
  NAND2_X1_LVT clock_module_0_i_36_10 (.ZN(clock_module_0_mclk_div_sel), .A1(
      clock_module_0_n_36_9), .A2(clock_module_0_n_36_1));
  AND2_X1_LVT clock_module_0_i_38_0 (.ZN(clock_module_0_mclk_div_en), .A1(
      clock_module_0_mclk_active), .A2(clock_module_0_mclk_div_sel));
  OR2_X1_LVT clock_module_0_clock_gate_mclk_i_0_0 (.ZN(
      clock_module_0_clock_gate_mclk_enable_in), .A1(clock_module_0_mclk_div_en), 
      .A2(scan_enable));
  INV_X1_LVT clock_module_0_clock_gate_mclk_i_1_0 (.ZN(
      clock_module_0_clock_gate_mclk_n_0), .A(dco_clk));
  DLH_X1_LVT clock_module_0_clock_gate_mclk_enable_latch_reg (.Q(
      clock_module_0_clock_gate_mclk_enable_latch), .D(
      clock_module_0_clock_gate_mclk_enable_in), .G(
      clock_module_0_clock_gate_mclk_n_0));
  AND2_X1_LVT clock_module_0_clock_gate_mclk_i_3_0 (.ZN(cpu_mclk), .A1(dco_clk), 
      .A2(clock_module_0_clock_gate_mclk_enable_latch));
  INV_X1_LVT clock_module_0_i_41_0 (.ZN(clock_module_0_dbg_rst_nxt), .A(dbg_en));
  INV_X1_LVT clock_module_0_sync_reset_por_i_0_0 (.ZN(
      clock_module_0_sync_reset_por_n_0), .A(clock_module_0_por_a));
  DFFS_X1_LVT \clock_module_0_sync_reset_por_data_sync_reg[0] (.Q(
      clock_module_0_sync_reset_por_n_1), .QN(), .CK(dco_clk), .D(1'b0), .SN(
      clock_module_0_sync_reset_por_n_0));
  DFFS_X1_LVT \clock_module_0_sync_reset_por_data_sync_reg[1] (.Q(
      clock_module_0_por_noscan), .QN(), .CK(dco_clk), .D(
      clock_module_0_sync_reset_por_n_1), .SN(clock_module_0_sync_reset_por_n_0));
  INV_X1_LVT clock_module_0_scan_mux_por_i_0_0 (.ZN(
      clock_module_0_scan_mux_por_n_0_0), .A(scan_mode));
  AOI22_X1_LVT clock_module_0_scan_mux_por_i_0_1 (.ZN(
      clock_module_0_scan_mux_por_n_0_1), .A1(clock_module_0_scan_mux_por_n_0_0), 
      .A2(clock_module_0_por_noscan), .B1(clock_module_0_por_a), .B2(scan_mode));
  INV_X1_LVT clock_module_0_scan_mux_por_i_0_2 (.ZN(por), .A(
      clock_module_0_scan_mux_por_n_0_1));
  INV_X1_LVT clock_module_0_i_3_0 (.ZN(clock_module_0_n_1), .A(por));
  DFFS_X1_LVT clock_module_0_dbg_rst_noscan_reg (.Q(
      clock_module_0_dbg_rst_noscan), .QN(), .CK(cpu_mclk), .D(
      clock_module_0_dbg_rst_nxt), .SN(clock_module_0_n_1));
  AND3_X1_LVT clock_module_0_i_46_0 (.ZN(clock_module_0_n_46_0), .A1(dbg_en), 
      .A2(puc_pnd_set), .A3(clock_module_0_dbg_rst_noscan));
  NOR2_X1_LVT clock_module_0_i_46_1 (.ZN(clock_module_0_n_28), .A1(
      clock_module_0_n_46_0), .A2(dbg_cpu_reset));
  OR2_X1_LVT clock_module_0_i_59_0 (.ZN(clock_module_0_puc_a), .A1(por), .A2(
      wdt_reset));
  INV_X1_LVT clock_module_0_scan_mux_puc_rst_a_i_0_0 (.ZN(
      clock_module_0_scan_mux_puc_rst_a_n_0_0), .A(scan_mode));
  AOI22_X1_LVT clock_module_0_scan_mux_puc_rst_a_i_0_1 (.ZN(
      clock_module_0_scan_mux_puc_rst_a_n_0_1), .A1(
      clock_module_0_scan_mux_puc_rst_a_n_0_0), .A2(clock_module_0_puc_a), .B1(
      clock_module_0_por_a), .B2(scan_mode));
  INV_X1_LVT clock_module_0_scan_mux_puc_rst_a_i_0_2 (.ZN(
      clock_module_0_puc_a_scan), .A(clock_module_0_scan_mux_puc_rst_a_n_0_1));
  INV_X1_LVT clock_module_0_sync_cell_puc_i_0_0 (.ZN(
      clock_module_0_sync_cell_puc_n_0), .A(clock_module_0_puc_a_scan));
  DFFR_X1_LVT \clock_module_0_sync_cell_puc_data_sync_reg[0] (.Q(
      clock_module_0_sync_cell_puc_n_1), .QN(), .CK(cpu_mclk), .D(
      clock_module_0_n_28), .RN(clock_module_0_sync_cell_puc_n_0));
  DFFR_X1_LVT \clock_module_0_sync_cell_puc_data_sync_reg[1] (.Q(
      clock_module_0_puc_noscan_n), .QN(), .CK(cpu_mclk), .D(
      clock_module_0_sync_cell_puc_n_1), .RN(clock_module_0_sync_cell_puc_n_0));
  INV_X1_LVT clock_module_0_i_21_0 (.ZN(puc_pnd_set), .A(
      clock_module_0_puc_noscan_n));
  INV_X1_LVT clock_module_0_scan_mux_puc_rst_i_0_0 (.ZN(
      clock_module_0_scan_mux_puc_rst_n_0_0), .A(scan_mode));
  AOI22_X1_LVT clock_module_0_scan_mux_puc_rst_i_0_1 (.ZN(
      clock_module_0_scan_mux_puc_rst_n_0_1), .A1(
      clock_module_0_scan_mux_puc_rst_n_0_0), .A2(puc_pnd_set), .B1(
      clock_module_0_por_a), .B2(scan_mode));
  INV_X1_LVT clock_module_0_scan_mux_puc_rst_i_0_2 (.ZN(puc_rst), .A(
      clock_module_0_scan_mux_puc_rst_n_0_1));
  INV_X1_LVT clock_module_0_i_18_0 (.ZN(clock_module_0_n_10), .A(puc_rst));
  DFFR_X1_LVT \clock_module_0_bcsctl1_reg[0] (.Q(clock_module_0_bcsctl1[0]), .QN(), 
      .CK(clock_module_0_n_9), .D(per_din[8]), .RN(clock_module_0_n_10));
  AND2_X1_LVT clock_module_0_and_cpuoff_mclk_dma_en_i_0_0 (.ZN(
      clock_module_0_cpuoff_and_mclk_dma_enable), .A1(clock_module_0_bcsctl1[0]), 
      .A2(mclk_dma_enable));
  AND2_X1_LVT clock_module_0_and_cpuoff_mclk_dma_wkup_i_0_0 (.ZN(
      clock_module_0_cpuoff_and_mclk_dma_wkup), .A1(clock_module_0_bcsctl1[0]), 
      .A2(mclk_dma_wkup));
  INV_X1_LVT clock_module_0_sync_cell_mclk_dma_wkup_i_0_0 (.ZN(
      clock_module_0_sync_cell_mclk_dma_wkup_n_0), .A(puc_rst));
  DFFR_X1_LVT \clock_module_0_sync_cell_mclk_dma_wkup_data_sync_reg[0] (.Q(
      clock_module_0_sync_cell_mclk_dma_wkup_n_1), .QN(), .CK(dco_clk), .D(
      clock_module_0_cpuoff_and_mclk_dma_wkup), .RN(
      clock_module_0_sync_cell_mclk_dma_wkup_n_0));
  DFFR_X1_LVT \clock_module_0_sync_cell_mclk_dma_wkup_data_sync_reg[1] (.Q(
      clock_module_0_cpuoff_and_mclk_dma_wkup_s), .QN(), .CK(dco_clk), .D(
      clock_module_0_sync_cell_mclk_dma_wkup_n_1), .RN(
      clock_module_0_sync_cell_mclk_dma_wkup_n_0));
  OR3_X1_LVT clock_module_0_i_39_0 (.ZN(clock_module_0_n_39_0), .A1(
      clock_module_0_cpuoff_and_mclk_dma_enable), .A2(clock_module_0_mclk_active), 
      .A3(clock_module_0_cpuoff_and_mclk_dma_wkup_s));
  AND2_X1_LVT clock_module_0_i_39_1 (.ZN(clock_module_0_mclk_dma_div_en), .A1(
      clock_module_0_n_39_0), .A2(clock_module_0_mclk_div_sel));
  OR2_X1_LVT clock_module_0_clock_gate_dma_mclk_i_0_0 (.ZN(
      clock_module_0_clock_gate_dma_mclk_enable_in), .A1(
      clock_module_0_mclk_dma_div_en), .A2(scan_enable));
  INV_X1_LVT clock_module_0_clock_gate_dma_mclk_i_1_0 (.ZN(
      clock_module_0_clock_gate_dma_mclk_n_0), .A(dco_clk));
  DLH_X1_LVT clock_module_0_clock_gate_dma_mclk_enable_latch_reg (.Q(
      clock_module_0_clock_gate_dma_mclk_enable_latch), .D(
      clock_module_0_clock_gate_dma_mclk_enable_in), .G(
      clock_module_0_clock_gate_dma_mclk_n_0));
  AND2_X1_LVT clock_module_0_clock_gate_dma_mclk_i_3_0 (.ZN(mclk), .A1(dco_clk), 
      .A2(clock_module_0_clock_gate_dma_mclk_enable_latch));
  CLKGATETST_X1_LVT clock_module_0_clk_gate_bcsctl1_reg (.GCK(clock_module_0_n_9), 
      .CK(mclk), .E(clock_module_0_bcsctl1_wr), .SE(1'b0));
  DFFR_X1_LVT \clock_module_0_bcsctl1_reg[5] (.Q(clock_module_0_bcsctl1[5]), .QN(), 
      .CK(clock_module_0_n_9), .D(per_din[13]), .RN(clock_module_0_n_10));
  INV_X1_LVT clock_module_0_i_28_2 (.ZN(clock_module_0_n_28_2), .A(
      clock_module_0_bcsctl1[5]));
  DFFR_X1_LVT \clock_module_0_bcsctl1_reg[4] (.Q(clock_module_0_bcsctl1[4]), .QN(), 
      .CK(clock_module_0_n_9), .D(per_din[12]), .RN(clock_module_0_n_10));
  OR2_X1_LVT clock_module_0_i_28_3 (.ZN(clock_module_0_n_28_3), .A1(
      clock_module_0_n_28_2), .A2(clock_module_0_bcsctl1[4]));
  INV_X1_LVT clock_module_0_i_23_0 (.ZN(clock_module_0_n_12), .A(
      clock_module_0_aclk_div[0]));
  OR2_X1_LVT clock_module_0_i_24_0 (.ZN(clock_module_0_n_15), .A1(
      clock_module_0_bcsctl1[4]), .A2(clock_module_0_bcsctl1[5]));
  CLKGATETST_X1_LVT clock_module_0_clk_gate_aclk_div_reg (.GCK(
      clock_module_0_n_11), .CK(dco_clk), .E(clock_module_0_n_15), .SE(1'b0));
  DFFR_X1_LVT \clock_module_0_aclk_div_reg[0] (.Q(clock_module_0_aclk_div[0]), 
      .QN(), .CK(clock_module_0_n_11), .D(clock_module_0_n_12), .RN(
      clock_module_0_n_10));
  HA_X1_LVT clock_module_0_i_23_1 (.CO(clock_module_0_n_23_0), .S(
      clock_module_0_n_13), .A(clock_module_0_aclk_div[1]), .B(
      clock_module_0_aclk_div[0]));
  DFFR_X1_LVT \clock_module_0_aclk_div_reg[1] (.Q(clock_module_0_aclk_div[1]), 
      .QN(), .CK(clock_module_0_n_11), .D(clock_module_0_n_13), .RN(
      clock_module_0_n_10));
  XNOR2_X1_LVT clock_module_0_i_23_2 (.ZN(clock_module_0_n_23_1), .A(
      clock_module_0_aclk_div[2]), .B(clock_module_0_n_23_0));
  INV_X1_LVT clock_module_0_i_23_3 (.ZN(clock_module_0_n_14), .A(
      clock_module_0_n_23_1));
  DFFR_X1_LVT \clock_module_0_aclk_div_reg[2] (.Q(clock_module_0_aclk_div[2]), 
      .QN(), .CK(clock_module_0_n_11), .D(clock_module_0_n_14), .RN(
      clock_module_0_n_10));
  AND3_X1_LVT clock_module_0_i_26_0 (.ZN(clock_module_0_n_16), .A1(
      clock_module_0_aclk_div[0]), .A2(clock_module_0_aclk_div[1]), .A3(
      clock_module_0_aclk_div[2]));
  INV_X1_LVT clock_module_0_i_28_4 (.ZN(clock_module_0_n_28_4), .A(
      clock_module_0_n_28_3));
  AND2_X1_LVT clock_module_0_i_27_0 (.ZN(clock_module_0_n_17), .A1(
      clock_module_0_aclk_div[0]), .A2(clock_module_0_aclk_div[1]));
  AOI22_X1_LVT clock_module_0_i_28_5 (.ZN(clock_module_0_n_28_5), .A1(
      clock_module_0_n_28_3), .A2(clock_module_0_n_16), .B1(
      clock_module_0_n_28_4), .B2(clock_module_0_n_17));
  INV_X1_LVT clock_module_0_i_28_6 (.ZN(clock_module_0_n_28_6), .A(
      clock_module_0_n_28_5));
  NAND2_X1_LVT clock_module_0_i_28_7 (.ZN(clock_module_0_n_28_7), .A1(
      clock_module_0_n_28_2), .A2(clock_module_0_bcsctl1[4]));
  INV_X1_LVT clock_module_0_i_28_8 (.ZN(clock_module_0_n_28_8), .A(
      clock_module_0_n_28_7));
  AOI22_X1_LVT clock_module_0_i_28_9 (.ZN(clock_module_0_n_28_9), .A1(
      clock_module_0_n_28_6), .A2(clock_module_0_n_28_7), .B1(
      clock_module_0_n_28_8), .B2(clock_module_0_aclk_div[0]));
  NOR2_X1_LVT clock_module_0_i_28_0 (.ZN(clock_module_0_n_28_0), .A1(
      clock_module_0_bcsctl1[4]), .A2(clock_module_0_bcsctl1[5]));
  INV_X1_LVT clock_module_0_i_28_1 (.ZN(clock_module_0_n_28_1), .A(
      clock_module_0_n_28_0));
  NAND2_X1_LVT clock_module_0_i_28_10 (.ZN(clock_module_0_aclk_div_sel), .A1(
      clock_module_0_n_28_9), .A2(clock_module_0_n_28_1));
  NAND2_X1_LVT clock_module_0_i_29_0 (.ZN(clock_module_0_n_29_0), .A1(cpu_en), 
      .A2(clock_module_0_aclk_div_sel));
  NOR2_X1_LVT clock_module_0_i_29_1 (.ZN(clock_module_0_aclk_div_en), .A1(
      clock_module_0_n_29_0), .A2(oscoff));
  OR2_X1_LVT clock_module_0_clock_gate_aclk_i_0_0 (.ZN(
      clock_module_0_clock_gate_aclk_enable_in), .A1(clock_module_0_aclk_div_en), 
      .A2(scan_enable));
  INV_X1_LVT clock_module_0_clock_gate_aclk_i_1_0 (.ZN(
      clock_module_0_clock_gate_aclk_n_0), .A(dco_clk));
  DLH_X1_LVT clock_module_0_clock_gate_aclk_enable_latch_reg (.Q(
      clock_module_0_clock_gate_aclk_enable_latch), .D(
      clock_module_0_clock_gate_aclk_enable_in), .G(
      clock_module_0_clock_gate_aclk_n_0));
  AND2_X1_LVT clock_module_0_clock_gate_aclk_i_3_0 (.ZN(aclk), .A1(dco_clk), .A2(
      clock_module_0_clock_gate_aclk_enable_latch));
  OR2_X1_LVT clock_module_0_clock_gate_dbg_clk_i_0_0 (.ZN(
      clock_module_0_clock_gate_dbg_clk_enable_in), .A1(dbg_en), .A2(scan_enable));
  INV_X1_LVT clock_module_0_clock_gate_dbg_clk_i_1_0 (.ZN(
      clock_module_0_clock_gate_dbg_clk_n_0), .A(cpu_mclk));
  DLH_X1_LVT clock_module_0_clock_gate_dbg_clk_enable_latch_reg (.Q(
      clock_module_0_clock_gate_dbg_clk_enable_latch), .D(
      clock_module_0_clock_gate_dbg_clk_enable_in), .G(
      clock_module_0_clock_gate_dbg_clk_n_0));
  AND2_X1_LVT clock_module_0_clock_gate_dbg_clk_i_3_0 (.ZN(dbg_clk), .A1(
      cpu_mclk), .A2(clock_module_0_clock_gate_dbg_clk_enable_latch));
  INV_X1_LVT clock_module_0_scan_mux_dbg_rst_i_0_0 (.ZN(
      clock_module_0_scan_mux_dbg_rst_n_0_0), .A(scan_mode));
  AOI22_X1_LVT clock_module_0_scan_mux_dbg_rst_i_0_1 (.ZN(
      clock_module_0_scan_mux_dbg_rst_n_0_1), .A1(
      clock_module_0_scan_mux_dbg_rst_n_0_0), .A2(clock_module_0_dbg_rst_noscan), 
      .B1(clock_module_0_por_a), .B2(scan_mode));
  INV_X1_LVT clock_module_0_scan_mux_dbg_rst_i_0_2 (.ZN(dbg_rst), .A(
      clock_module_0_scan_mux_dbg_rst_n_0_1));
  DFFR_X1_LVT \clock_module_0_bcsctl2_reg[7] (.Q(clock_module_0_bcsctl2[7]), .QN(), 
      .CK(clock_module_0_n_8), .D(1'b0), .RN(clock_module_0_n_10));
  INV_X1_LVT clock_module_0_i_58_0 (.ZN(clock_module_0_n_39), .A(
      clock_module_0_bcsctl2[7]));
  AND2_X1_LVT clock_module_0_and_dco_mclk_wkup_i_0_0 (.ZN(
      clock_module_0_dco_mclk_wkup), .A1(mclk_wkup), .A2(clock_module_0_n_39));
  INV_X1_LVT clock_module_0_i_57_0 (.ZN(clock_module_0_n_38), .A(dco_enable));
  AND2_X1_LVT clock_module_0_and_cpuoff_mclk_en_i_0_0 (.ZN(
      clock_module_0_cpuoff_and_mclk_enable), .A1(cpuoff), .A2(mclk_enable));
  AND2_X1_LVT clock_module_0_and_dco_dis1_i_0_0 (.ZN(
      clock_module_0_cpu_enabled_with_dco), .A1(clock_module_0_n_39), .A2(
      clock_module_0_cpuoff_and_mclk_enable));
  DFFR_X1_LVT \clock_module_0_bcsctl1_reg[2] (.Q(clock_module_0_bcsctl1[2]), .QN(), 
      .CK(clock_module_0_n_9), .D(per_din[10]), .RN(clock_module_0_n_10));
  AND2_X1_LVT clock_module_0_and_scg0_mclk_dma_en_i_0_0 (.ZN(
      clock_module_0_scg0_and_mclk_dma_enable), .A1(clock_module_0_bcsctl1[2]), 
      .A2(mclk_dma_enable));
  NOR2_X1_LVT clock_module_0_i_60_0 (.ZN(clock_module_0_n_40), .A1(
      clock_module_0_cpu_enabled_with_dco), .A2(
      clock_module_0_scg0_and_mclk_dma_enable));
  AND2_X1_LVT clock_module_0_and_dco_dis2_i_0_0 (.ZN(
      clock_module_0_dco_not_enabled_by_dbg), .A1(clock_module_0_dbg_rst_nxt), 
      .A2(clock_module_0_n_40));
  AND2_X1_LVT clock_module_0_and_dco_dis3_i_0_0 (.ZN(
      clock_module_0_dco_disable_by_scg0), .A1(scg0), .A2(
      clock_module_0_dco_not_enabled_by_dbg));
  INV_X1_LVT clock_module_0_i_42_0 (.ZN(clock_module_0_n_25), .A(
      clock_module_0_dco_disable_by_scg0));
  INV_X1_LVT clock_module_0_i_55_0 (.ZN(clock_module_0_n_36), .A(cpu_en));
  INV_X1_LVT clock_module_0_i_56_0 (.ZN(clock_module_0_n_37), .A(mclk_enable));
  AND2_X1_LVT clock_module_0_and_dco_dis4_i_0_0 (.ZN(
      clock_module_0_dco_disable_by_cpu_en), .A1(clock_module_0_n_36), .A2(
      clock_module_0_n_37));
  INV_X1_LVT clock_module_0_i_43_0 (.ZN(clock_module_0_n_26), .A(
      clock_module_0_dco_disable_by_cpu_en));
  AND2_X1_LVT clock_module_0_and_dco_dis5_i_0_0 (.ZN(
      clock_module_0_dco_enable_nxt), .A1(clock_module_0_n_25), .A2(
      clock_module_0_n_26));
  AND2_X1_LVT clock_module_0_and_dco_en_wkup_i_0_0 (.ZN(
      clock_module_0_dco_en_wkup), .A1(clock_module_0_n_38), .A2(
      clock_module_0_dco_enable_nxt));
  AND2_X1_LVT clock_module_0_and_scg0_mclk_dma_wkup_i_0_0 (.ZN(
      clock_module_0_scg0_and_mclk_dma_wkup), .A1(clock_module_0_bcsctl1[2]), 
      .A2(mclk_dma_wkup));
  OR3_X1_LVT clock_module_0_i_44_0 (.ZN(clock_module_0_dco_wkup_set), .A1(
      clock_module_0_dco_mclk_wkup), .A2(clock_module_0_dco_en_wkup), .A3(
      clock_module_0_scg0_and_mclk_dma_wkup));
  INV_X1_LVT clock_module_0_scan_mux_dco_wkup_observe_i_0_0 (.ZN(
      clock_module_0_scan_mux_dco_wkup_observe_n_0_0), .A(scan_mode));
  AOI22_X1_LVT clock_module_0_scan_mux_dco_wkup_observe_i_0_1 (.ZN(
      clock_module_0_scan_mux_dco_wkup_observe_n_0_1), .A1(
      clock_module_0_scan_mux_dco_wkup_observe_n_0_0), .A2(1'b0), .B1(
      clock_module_0_dco_wkup_set), .B2(scan_mode));
  INV_X1_LVT clock_module_0_scan_mux_dco_wkup_observe_i_0_2 (.ZN(
      clock_module_0_dco_wkup_set_scan_observe), .A(
      clock_module_0_scan_mux_dco_wkup_observe_n_0_1));
  INV_X1_LVT clock_module_0_i_1_0 (.ZN(clock_module_0_n_1_0), .A(
      clock_module_0_dco_wkup_set_scan_observe));
  NAND2_X1_LVT clock_module_0_i_1_1 (.ZN(clock_module_0_n_0), .A1(
      clock_module_0_n_1_0), .A2(clock_module_0_dco_enable_nxt));
  DFFS_X1_LVT clock_module_0_dco_disable_reg (.Q(clock_module_0_dco_disable), 
      .QN(), .CK(dco_clk), .D(clock_module_0_n_0), .SN(clock_module_0_n_1));
  INV_X1_LVT clock_module_0_i_5_0 (.ZN(clock_module_0_n_2), .A(
      clock_module_0_dco_disable));
  INV_X1_LVT clock_module_0_i_0_0 (.ZN(clock_module_0_nodiv_mclk_n), .A(dco_clk));
  DFFR_X1_LVT clock_module_0_dco_enable_reg (.Q(dco_enable), .QN(), .CK(
      clock_module_0_nodiv_mclk_n), .D(clock_module_0_n_2), .RN(
      clock_module_0_n_1));
  OR2_X1_LVT clock_module_0_i_61_0 (.ZN(clock_module_0_n_41), .A1(
      clock_module_0_dco_wkup_set), .A2(por));
  INV_X1_LVT clock_module_0_scan_mux_dco_wkup_i_0_0 (.ZN(
      clock_module_0_scan_mux_dco_wkup_n_0_0), .A(scan_mode));
  AOI22_X1_LVT clock_module_0_scan_mux_dco_wkup_i_0_1 (.ZN(
      clock_module_0_scan_mux_dco_wkup_n_0_1), .A1(
      clock_module_0_scan_mux_dco_wkup_n_0_0), .A2(clock_module_0_n_41), .B1(
      clock_module_0_por_a), .B2(scan_mode));
  INV_X1_LVT clock_module_0_scan_mux_dco_wkup_i_0_2 (.ZN(
      clock_module_0_dco_wkup_set_scan), .A(
      clock_module_0_scan_mux_dco_wkup_n_0_1));
  INV_X1_LVT clock_module_0_sync_cell_dco_wkup_i_0_0 (.ZN(
      clock_module_0_sync_cell_dco_wkup_n_0), .A(
      clock_module_0_dco_wkup_set_scan));
  DFFR_X1_LVT \clock_module_0_sync_cell_dco_wkup_data_sync_reg[0] (.Q(
      clock_module_0_sync_cell_dco_wkup_n_1), .QN(), .CK(
      clock_module_0_nodiv_mclk_n), .D(1'b1), .RN(
      clock_module_0_sync_cell_dco_wkup_n_0));
  DFFR_X1_LVT \clock_module_0_sync_cell_dco_wkup_data_sync_reg[1] (.Q(
      clock_module_0_dco_wkup_n), .QN(), .CK(clock_module_0_nodiv_mclk_n), .D(
      clock_module_0_sync_cell_dco_wkup_n_1), .RN(
      clock_module_0_sync_cell_dco_wkup_n_0));
  INV_X1_LVT clock_module_0_i_45_0 (.ZN(clock_module_0_n_27), .A(
      clock_module_0_dco_wkup_n));
  AND2_X1_LVT clock_module_0_and_dco_wkup_i_0_0 (.ZN(dco_wkup), .A1(
      clock_module_0_n_27), .A2(cpu_en));
  NOR2_X1_LVT clock_module_0_i_8_0 (.ZN(clock_module_0_n_3), .A1(per_we[0]), .A2(
      per_we[1]));
  AND2_X1_LVT clock_module_0_i_9_0 (.ZN(clock_module_0_reg_read), .A1(
      clock_module_0_n_3), .A2(clock_module_0_reg_sel));
  AND2_X1_LVT clock_module_0_i_12_0 (.ZN(clock_module_0_n_6), .A1(
      clock_module_0_reg_read), .A2(clock_module_0_n_5));
  DFFR_X1_LVT \clock_module_0_bcsctl1_reg[7] (.Q(clock_module_0_bcsctl1[7]), .QN(), 
      .CK(clock_module_0_n_9), .D(1'b0), .RN(clock_module_0_n_10));
  AND2_X1_LVT clock_module_0_i_20_15 (.ZN(per_dout_clk[15]), .A1(
      clock_module_0_n_6), .A2(clock_module_0_bcsctl1[7]));
  DFFR_X1_LVT \clock_module_0_bcsctl1_reg[6] (.Q(clock_module_0_bcsctl1[6]), .QN(), 
      .CK(clock_module_0_n_9), .D(1'b0), .RN(clock_module_0_n_10));
  AND2_X1_LVT clock_module_0_i_20_14 (.ZN(per_dout_clk[14]), .A1(
      clock_module_0_n_6), .A2(clock_module_0_bcsctl1[6]));
  AND2_X1_LVT clock_module_0_i_20_13 (.ZN(per_dout_clk[13]), .A1(
      clock_module_0_n_6), .A2(clock_module_0_bcsctl1[5]));
  AND2_X1_LVT clock_module_0_i_20_12 (.ZN(per_dout_clk[12]), .A1(
      clock_module_0_n_6), .A2(clock_module_0_bcsctl1[4]));
  DFFR_X1_LVT \clock_module_0_bcsctl1_reg[3] (.Q(clock_module_0_bcsctl1[3]), .QN(), 
      .CK(clock_module_0_n_9), .D(per_din[11]), .RN(clock_module_0_n_10));
  AND2_X1_LVT clock_module_0_i_20_11 (.ZN(per_dout_clk[11]), .A1(
      clock_module_0_n_6), .A2(clock_module_0_bcsctl1[3]));
  AND2_X1_LVT clock_module_0_i_20_10 (.ZN(per_dout_clk[10]), .A1(
      clock_module_0_n_6), .A2(clock_module_0_bcsctl1[2]));
  DFFR_X1_LVT \clock_module_0_bcsctl1_reg[1] (.Q(clock_module_0_bcsctl1[1]), .QN(), 
      .CK(clock_module_0_n_9), .D(1'b0), .RN(clock_module_0_n_10));
  AND2_X1_LVT clock_module_0_i_20_9 (.ZN(per_dout_clk[9]), .A1(
      clock_module_0_n_6), .A2(clock_module_0_bcsctl1[1]));
  AND2_X1_LVT clock_module_0_i_20_8 (.ZN(per_dout_clk[8]), .A1(
      clock_module_0_bcsctl1[0]), .A2(clock_module_0_n_6));
  AND2_X1_LVT clock_module_0_i_12_1 (.ZN(clock_module_0_n_7), .A1(
      clock_module_0_reg_read), .A2(clock_module_0_n_4));
  AND2_X1_LVT clock_module_0_i_20_7 (.ZN(per_dout_clk[7]), .A1(
      clock_module_0_n_7), .A2(clock_module_0_bcsctl2[7]));
  DFFR_X1_LVT \clock_module_0_bcsctl2_reg[6] (.Q(clock_module_0_bcsctl2[6]), .QN(), 
      .CK(clock_module_0_n_8), .D(1'b0), .RN(clock_module_0_n_10));
  AND2_X1_LVT clock_module_0_i_20_6 (.ZN(per_dout_clk[6]), .A1(
      clock_module_0_n_7), .A2(clock_module_0_bcsctl2[6]));
  AND2_X1_LVT clock_module_0_i_20_5 (.ZN(per_dout_clk[5]), .A1(
      clock_module_0_n_7), .A2(clock_module_0_bcsctl2[5]));
  AND2_X1_LVT clock_module_0_i_20_4 (.ZN(per_dout_clk[4]), .A1(
      clock_module_0_n_7), .A2(clock_module_0_bcsctl2[4]));
  DFFR_X1_LVT \clock_module_0_bcsctl2_reg[3] (.Q(clock_module_0_bcsctl2[3]), .QN(), 
      .CK(clock_module_0_n_8), .D(1'b0), .RN(clock_module_0_n_10));
  AND2_X1_LVT clock_module_0_i_20_3 (.ZN(per_dout_clk[3]), .A1(
      clock_module_0_n_7), .A2(clock_module_0_bcsctl2[3]));
  DFFR_X1_LVT \clock_module_0_bcsctl2_reg[2] (.Q(clock_module_0_bcsctl2[2]), .QN(), 
      .CK(clock_module_0_n_8), .D(per_din[2]), .RN(clock_module_0_n_10));
  AND2_X1_LVT clock_module_0_i_20_2 (.ZN(per_dout_clk[2]), .A1(
      clock_module_0_n_7), .A2(clock_module_0_bcsctl2[2]));
  DFFR_X1_LVT \clock_module_0_bcsctl2_reg[1] (.Q(clock_module_0_bcsctl2[1]), .QN(), 
      .CK(clock_module_0_n_8), .D(per_din[1]), .RN(clock_module_0_n_10));
  AND2_X1_LVT clock_module_0_i_20_1 (.ZN(per_dout_clk[1]), .A1(
      clock_module_0_n_7), .A2(clock_module_0_bcsctl2[1]));
  DFFR_X1_LVT \clock_module_0_bcsctl2_reg[0] (.Q(clock_module_0_bcsctl2[0]), .QN(), 
      .CK(clock_module_0_n_8), .D(1'b0), .RN(clock_module_0_n_10));
  AND2_X1_LVT clock_module_0_i_20_0 (.ZN(per_dout_clk[0]), .A1(
      clock_module_0_bcsctl2[0]), .A2(clock_module_0_n_7));
  INV_X1_LVT clock_module_0_i_54_0 (.ZN(clock_module_0_n_54_0), .A(scg1));
  AND2_X1_LVT clock_module_0_and_scg1_mclk_dma_wkup_i_0_0 (.ZN(
      clock_module_0_scg1_and_mclk_dma_wkup), .A1(clock_module_0_bcsctl1[3]), 
      .A2(mclk_dma_wkup));
  INV_X1_LVT clock_module_0_sync_cell_smclk_dma_wkup_i_0_0 (.ZN(
      clock_module_0_sync_cell_smclk_dma_wkup_n_0), .A(puc_rst));
  DFFR_X1_LVT \clock_module_0_sync_cell_smclk_dma_wkup_data_sync_reg[0] (.Q(
      clock_module_0_sync_cell_smclk_dma_wkup_n_1), .QN(), .CK(dco_clk), .D(
      clock_module_0_scg1_and_mclk_dma_wkup), .RN(
      clock_module_0_sync_cell_smclk_dma_wkup_n_0));
  DFFR_X1_LVT \clock_module_0_sync_cell_smclk_dma_wkup_data_sync_reg[1] (.Q(
      clock_module_0_scg1_and_mclk_dma_wkup_s), .QN(), .CK(dco_clk), .D(
      clock_module_0_sync_cell_smclk_dma_wkup_n_1), .RN(
      clock_module_0_sync_cell_smclk_dma_wkup_n_0));
  AND2_X1_LVT clock_module_0_and_scg1_mclk_dma_en_i_0_0 (.ZN(
      clock_module_0_scg1_and_mclk_dma_enable), .A1(clock_module_0_bcsctl1[3]), 
      .A2(mclk_dma_enable));
  NOR3_X1_LVT clock_module_0_i_54_1 (.ZN(clock_module_0_n_54_1), .A1(
      clock_module_0_n_54_0), .A2(clock_module_0_scg1_and_mclk_dma_wkup_s), .A3(
      clock_module_0_scg1_and_mclk_dma_enable));
  INV_X1_LVT clock_module_0_i_53_2 (.ZN(clock_module_0_n_53_2), .A(
      clock_module_0_bcsctl2[2]));
  OR2_X1_LVT clock_module_0_i_53_3 (.ZN(clock_module_0_n_53_3), .A1(
      clock_module_0_n_53_2), .A2(clock_module_0_bcsctl2[1]));
  INV_X1_LVT clock_module_0_i_48_0 (.ZN(clock_module_0_n_30), .A(
      clock_module_0_smclk_div[0]));
  OR2_X1_LVT clock_module_0_i_49_0 (.ZN(clock_module_0_n_33), .A1(
      clock_module_0_bcsctl2[1]), .A2(clock_module_0_bcsctl2[2]));
  CLKGATETST_X1_LVT clock_module_0_clk_gate_smclk_div_reg (.GCK(
      clock_module_0_n_29), .CK(dco_clk), .E(clock_module_0_n_33), .SE(1'b0));
  DFFR_X1_LVT \clock_module_0_smclk_div_reg[0] (.Q(clock_module_0_smclk_div[0]), 
      .QN(), .CK(clock_module_0_n_29), .D(clock_module_0_n_30), .RN(
      clock_module_0_n_10));
  HA_X1_LVT clock_module_0_i_48_1 (.CO(clock_module_0_n_48_0), .S(
      clock_module_0_n_31), .A(clock_module_0_smclk_div[1]), .B(
      clock_module_0_smclk_div[0]));
  DFFR_X1_LVT \clock_module_0_smclk_div_reg[1] (.Q(clock_module_0_smclk_div[1]), 
      .QN(), .CK(clock_module_0_n_29), .D(clock_module_0_n_31), .RN(
      clock_module_0_n_10));
  XNOR2_X1_LVT clock_module_0_i_48_2 (.ZN(clock_module_0_n_48_1), .A(
      clock_module_0_smclk_div[2]), .B(clock_module_0_n_48_0));
  INV_X1_LVT clock_module_0_i_48_3 (.ZN(clock_module_0_n_32), .A(
      clock_module_0_n_48_1));
  DFFR_X1_LVT \clock_module_0_smclk_div_reg[2] (.Q(clock_module_0_smclk_div[2]), 
      .QN(), .CK(clock_module_0_n_29), .D(clock_module_0_n_32), .RN(
      clock_module_0_n_10));
  AND3_X1_LVT clock_module_0_i_51_0 (.ZN(clock_module_0_n_34), .A1(
      clock_module_0_smclk_div[0]), .A2(clock_module_0_smclk_div[1]), .A3(
      clock_module_0_smclk_div[2]));
  INV_X1_LVT clock_module_0_i_53_4 (.ZN(clock_module_0_n_53_4), .A(
      clock_module_0_n_53_3));
  AND2_X1_LVT clock_module_0_i_52_0 (.ZN(clock_module_0_n_35), .A1(
      clock_module_0_smclk_div[0]), .A2(clock_module_0_smclk_div[1]));
  AOI22_X1_LVT clock_module_0_i_53_5 (.ZN(clock_module_0_n_53_5), .A1(
      clock_module_0_n_53_3), .A2(clock_module_0_n_34), .B1(
      clock_module_0_n_53_4), .B2(clock_module_0_n_35));
  INV_X1_LVT clock_module_0_i_53_6 (.ZN(clock_module_0_n_53_6), .A(
      clock_module_0_n_53_5));
  NAND2_X1_LVT clock_module_0_i_53_7 (.ZN(clock_module_0_n_53_7), .A1(
      clock_module_0_n_53_2), .A2(clock_module_0_bcsctl2[1]));
  INV_X1_LVT clock_module_0_i_53_8 (.ZN(clock_module_0_n_53_8), .A(
      clock_module_0_n_53_7));
  AOI22_X1_LVT clock_module_0_i_53_9 (.ZN(clock_module_0_n_53_9), .A1(
      clock_module_0_n_53_6), .A2(clock_module_0_n_53_7), .B1(
      clock_module_0_n_53_8), .B2(clock_module_0_smclk_div[0]));
  NOR2_X1_LVT clock_module_0_i_53_0 (.ZN(clock_module_0_n_53_0), .A1(
      clock_module_0_bcsctl2[1]), .A2(clock_module_0_bcsctl2[2]));
  INV_X1_LVT clock_module_0_i_53_1 (.ZN(clock_module_0_n_53_1), .A(
      clock_module_0_n_53_0));
  NAND2_X1_LVT clock_module_0_i_53_10 (.ZN(clock_module_0_smclk_div_sel), .A1(
      clock_module_0_n_53_9), .A2(clock_module_0_n_53_1));
  NAND2_X1_LVT clock_module_0_i_54_2 (.ZN(clock_module_0_n_54_2), .A1(cpu_en), 
      .A2(clock_module_0_smclk_div_sel));
  NOR2_X1_LVT clock_module_0_i_54_3 (.ZN(clock_module_0_smclk_div_en), .A1(
      clock_module_0_n_54_1), .A2(clock_module_0_n_54_2));
  OR2_X1_LVT clock_module_0_clock_gate_smclk_i_0_0 (.ZN(
      clock_module_0_clock_gate_smclk_enable_in), .A1(
      clock_module_0_smclk_div_en), .A2(scan_enable));
  INV_X1_LVT clock_module_0_clock_gate_smclk_i_1_0 (.ZN(
      clock_module_0_clock_gate_smclk_n_0), .A(dco_clk));
  DLH_X1_LVT clock_module_0_clock_gate_smclk_enable_latch_reg (.Q(
      clock_module_0_clock_gate_smclk_enable_latch), .D(
      clock_module_0_clock_gate_smclk_enable_in), .G(
      clock_module_0_clock_gate_smclk_n_0));
  AND2_X1_LVT clock_module_0_clock_gate_smclk_i_3_0 (.ZN(smclk), .A1(dco_clk), 
      .A2(clock_module_0_clock_gate_smclk_enable_latch));
endmodule

