module has_bigger_constant_value(A,C);
   input [120:0]A;
   output [120:0]C;
   wire [63:0]slongv;
  assign slongv[63] = 1'b0;
  assign slongv[62] = 1'b0;
  assign slongv[61] = 1'b0;
  assign slongv[60] = 1'b0;
  assign slongv[59] = 1'b1;
  assign slongv[58] = 1'b0;
  assign slongv[57] = 1'b1;
  assign slongv[56] = 1'b1;
  assign slongv[55] = 1'b1;
  assign slongv[54] = 1'b1;
  assign slongv[53] = 1'b0;
  assign slongv[52] = 1'b1;
  assign slongv[51] = 1'bx;
  assign slongv[50] = 1'bz;
  assign slongv[49] = 1'bx;
  assign slongv[48] = 1'bz;
  assign slongv[47] = 1'bz;
  assign slongv[46] = 1'bx;
  assign slongv[45] = 1'bz;
  assign slongv[44] = 1'bx;
  assign slongv[43] = 1'bz;
  assign slongv[42] = 1'bz;
  assign slongv[41] = 1'bz;
  assign slongv[40] = 1'bz;
  assign slongv[39] = 1'bx;
  assign slongv[38] = 1'bx;
  assign slongv[37] = 1'bx;
  assign slongv[36] = 1'bx;
  assign slongv[35] = 1'b0;
  assign slongv[34] = 1'b0;
  assign slongv[33] = 1'b0;
  assign slongv[32] = 1'b0;
  assign slongv[31] = A[31];
  assign slongv[30] = A[30];
  assign slongv[29] = A[29];
  assign slongv[28] = A[28];
  assign slongv[27] = A[27];
  assign slongv[26] = A[26];
  assign slongv[25] = A[25];
  assign slongv[24] = A[24];
  assign slongv[23] = A[23];
  assign slongv[22] = A[22];
  assign slongv[21] = A[21];
  assign slongv[20] = A[20];
  assign slongv[19] = A[19];
  assign slongv[18] = A[18];
  assign slongv[17] = A[17];
  assign slongv[16] = A[16];
  assign slongv[15] = A[15];
  assign slongv[14] = A[14];
  assign slongv[13] = A[13];
  assign slongv[12] = A[12];
  assign slongv[11] = A[11];
  assign slongv[10] = A[10];
  assign slongv[9] = A[9];
  assign slongv[8] = A[8];
  assign slongv[7] = A[7];
  assign slongv[6] = A[6];
  assign slongv[5] = A[5];
  assign slongv[4] = A[4];
  assign slongv[3] = A[3];
  assign slongv[2] = A[2];
  assign slongv[1] = A[1];
  assign slongv[0] = A[0];
  assign C[120] = A[120];
  assign C[119] = A[119];
  assign C[118] = A[118];
  assign C[117] = A[117];
  assign C[116] = A[116];
  assign C[115] = A[115];
  assign C[114] = A[114];
  assign C[113] = A[113];
  assign C[112] = A[112];
  assign C[111] = A[111];
  assign C[110] = A[110];
  assign C[109] = A[109];
  assign C[108] = A[108];
  assign C[107] = A[107];
  assign C[106] = A[106];
  assign C[105] = A[105];
  assign C[104] = A[104];
  assign C[103] = A[103];
  assign C[102] = A[102];
  assign C[101] = A[101];
  assign C[100] = A[100];
  assign C[99] = A[99];
  assign C[98] = A[98];
  assign C[97] = A[97];
  assign C[96] = A[96];
  assign C[95] = A[95];
  assign C[94] = A[94];
  assign C[93] = A[93];
  assign C[92] = A[92];
  assign C[91] = A[91];
  assign C[90] = A[90];
  assign C[89] = A[89];
  assign C[88] = A[88];
  assign C[87] = A[87];
  assign C[86] = A[86];
  assign C[85] = A[85];
  assign C[84] = A[84];
  assign C[83] = A[83];
  assign C[82] = A[82];
  assign C[81] = A[81];
  assign C[80] = A[80];
  assign C[79] = A[79];
  assign C[78] = A[78];
  assign C[77] = A[77];
  assign C[76] = A[76];
  assign C[75] = A[75];
  assign C[74] = A[74];
  assign C[73] = A[73];
  assign C[72] = A[72];
  assign C[71] = A[71];
  assign C[70] = A[70];
  assign C[69] = A[69];
  assign C[68] = A[68];
  assign C[67] = A[67];
  assign C[66] = A[66];
  assign C[65] = A[65];
  assign C[64] = A[64];
  assign C[63] = A[63];
  assign C[62] = A[62];
  assign C[61] = A[61];
  assign C[60] = A[60];
  assign C[59] = A[59];
  assign C[58] = A[58];
  assign C[57] = A[57];
  assign C[56] = A[56];
  assign C[55] = A[55];
  assign C[54] = A[54];
  assign C[53] = A[53];
  assign C[52] = A[52];
  assign C[51] = A[51];
  assign C[50] = A[50];
  assign C[49] = A[49];
  assign C[48] = A[48];
  assign C[47] = A[47];
  assign C[46] = A[46];
  assign C[45] = A[45];
  assign C[44] = A[44];
  assign C[43] = A[43];
  assign C[42] = A[42];
  assign C[41] = A[41];
  assign C[40] = A[40];
  assign C[39] = A[39];
  assign C[38] = A[38];
  assign C[37] = A[37];
  assign C[36] = A[36];
  assign C[35] = A[35];
  assign C[34] = A[34];
  assign C[33] = A[33];
  assign C[32] = A[32];
  assign C[31] = A[31];
  assign C[30] = A[30];
  assign C[29] = A[29];
  assign C[28] = A[28];
  assign C[27] = A[27];
  assign C[26] = A[26];
  assign C[25] = A[25];
  assign C[24] = A[24];
  assign C[23] = A[23];
  assign C[22] = A[22];
  assign C[21] = A[21];
  assign C[20] = A[20];
  assign C[19] = A[19];
  assign C[18] = A[18];
  assign C[17] = A[17];
  assign C[16] = A[16];
  assign C[15] = A[15];
  assign C[14] = A[14];
  assign C[13] = A[13];
  assign C[12] = A[12];
  assign C[11] = A[11];
  assign C[10] = A[10];
  assign C[9] = A[9];
  assign C[8] = A[8];
  assign C[7] = A[7];
  assign C[6] = A[6];
  assign C[5] = A[5];
  assign C[4] = A[4];
  assign C[3] = A[3];
  assign C[2] = A[2];
  assign C[1] = A[1];
  assign C[0] = A[0];
endmodule

